MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       8bz�|�|�|�u{��n�u{���[�o�y�|�&�u{��U�u{��}�u{��}�Rich|�                PE  L ��R        � "!	  �   n      �      �                          P                              ��  N   ��  <                            0 �
  p�                             �  @            �  4                          .text   ز      �                    `.rdata  �)   �   *   �              @  @.data   �,         �              @  �.reloc  &   0     �              @  B                                                                                                                                                                                                                                                                                                                                                                                                        U��E��u�E�M�h�d�   ]� �����������U����  � 3ŉE��=l �  VWh  �8  ����hh  VP�� j\V�%  ��+��OQ������VR��  ��������Ƅ=���� H�H@��u��@� �D� �f�H� �P������Rf�H��  V��  ������h<� P�  ������u>Ph$� h� �,� P�(� h�� �  ��_^�M�3��  ��]����$    W�����h�  Q�>  j�����h�� R���i  ����t��u��33����$    ������������@��u퍅����Ph�� �  ��W�  ��������O�GG��u�f��� ������f�H�H@��u���� ��� ���� �H�P������H��$    �H@��u���� ��� �j�Pj ������P� � �l��u/�5,� Ph$� h�� �֋=(� P��j h$� ������Q��P��_^�M�3��F  ��]���������������U�������lhL� P�� ��t]��3�]Ë�U��]��  �U��W�}3�������ك��E���8t3�����_�Ë�U��SV�uW3����;�u�v  WWWWW�    ��  ����B�F�t7V�!  V����
  V�
  P��	  ����}�����F;�t
P�  Y�~�~��_^[]�jh�� �  �M��3��u3�;���;�u��  �    WWWWW�{  �������F@t�~�E��  �V��  Y�}�V�*���Y�E��E������   �ՋuV�1  YË�U��Q�e� S�]��u3��   W��ru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+���jh�� ��  �E�E��E�3�;�u$9]t�  �    SSSSS�?  ��3���   3�9]��;�t�3��u;���;�t�9]tډu�V�  Y�]��F@uvV��  Y���t���t�����ȃ�������H�A$u)���t���t������������H�@$�t�  �    SSSSS�  ���]�9]�t<�}��Mt2�Nx
��A��V��  Y�E؃��u
;}u�]���G�}�<
uɈ�E������   �E���  Ëu�V�)  Y�jh � �  3ۉ]�3��};���;�u�p  �    SSSSS��
  ��3��y3��u;���;�t�3�8��;�t���  �E;�u�/  �    �ʉ]�8u �  �    j��E�Ph ��  ���P�uVW�  ���E��E������	   �E��   ��u�e  YË�U��j@�u�u�*�����]Ë�U��]�"  jh � �  3�3�9u��;�u�
  �    VVVVV�
  ������_�
  j [�Pj��  YY�u��
  �P�f  Y���EPV�u�
  �P�K  �E��|
  �PW��  ���E������	   �E��X  ��V
  �� Pj��  YYá ��3�9p�����������������̋L$W����   VS�ًt$��   �|$u����   �'��������t+��t/��   u����ua��t��������t7��u�D$[^_���   t�������   ��   u����ut�����u�[^�D$_É����t�����~�Ѓ��3��� �t܄�t,��t��  � t��   �uĉ�����  �����   ��3҉��3���t3������u����w����D$[^_�; u���Q#  ��U��EVW��u|P��2  Y��u3��  �(  ��u�3  ���2  �� ��,�A1  �x�t  ��}�(%  ���l0  ��| ��-  ��|j �+  Y��u�t�   �  ��3�;�u19=t~��t9=u�K-  9}u{�b  ��$  �z2  �j��uY�$  h  j��)  ��YY;��6���V�5��5���#  Y�Ѕ�tWV�$  YY�� �N���V�  Y�������uW�<'  Y3�@_^]� jh@� �h	  ����]3�@�E��u9t��   �e� ;�t��u.�X� ��tWVS�ЉE�}� ��   WVS�r����E����   WVS�����E��u$��u WPS����Wj S�B����X� ��tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�X� ��tWVS�ЉE��E������E���E��	PQ��2  YYËe��E�����3���  Ë�U��}u��2  �u�M�U�����Y]� ��Vjh ���f3  �`� ��^��`� ��3  ��U��V���`� �3  �EtV�]���Y��^]� ��U��V�u���73  �`� ��^]� ��U�����u�P6  Y��t�u�j5  Y��t�������u�����T���h�� ��4  YV�M�����h\� �E�P�&6  �jh�� �  �u��tu�=PuCj��7  Y�e� V��7  Y�E��t	VP�8  YY�E������   �}� u7�u�
j�6  Y�Vj �5$�� ��u�  ���� P��  �Y�D  Ë�U��V�uWV�MC  Y���tP����u	���   u��u�@Dtj�"C  j���C  YY;�tV�C  YP�� ��u
�� ���3�V�iB  �����������Y�D0 ��tW�  Y����3�_^]�jh�� �V  �E���u�\  �  �A  � 	   ����   3�;�|;lr!�3  �8�  � 	   WWWWW�  ���ɋ��������������L1��t�P�B  Y�}���D0t�u�����Y�E���  � 	   �M���E������	   �E���  ��u�C  YË�U��EV3�;�u�  VVVVV�    �	  �������@^]Ë�U��V�u�F��t�t�v�����f����3�Y��F�F^]Ë�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�i���YP�aK  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV� ���P��K  Y��Y��3�^]�jh�� �v  3��}�}�j��4  Y�}�3��u�;5�,��   ����98t^� �@�tVPV�  YY3�B�U������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��uࡄ�4�V�  YY��E������   �}�E�t�E���  �j�13  Y�j����YË�U��E��]Ë�U���(  � 3ŉE������� SjL������j P�K  ��������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������0� j ���,� ��(���P�(� ��u��uj�J  Yh ��$� P� � �M�3�[�����Ë�U���5��  Y��t]��j�pJ  Y]������U��E3�;�X tA��-r�H��wjX]Ë�\ ]�D���jY;��#���]���  ��u��Ã����  ��u��Ã�Ë�U��V������MQ�����Y�������0^]ø�á�,Vj^��u�   �;�}�ƣ�,jP�!  YY����ujV�5�,�o!  YY����ujX^�3ҹ������� ����H|�j�^3ҹ�W�����������������t;�t��u�1�� B��8|�_3�^��S����= t�I  �5��V���YË�U��V�u��;�r"��(w��+�����Q�1  �N �  Y�
�� V�4� ^]Ë�U��E��}��P��0  �E�H �  Y]ËE�� P�4� ]Ë�U��E��;�r=(w�`���+�����P��/  Y]Ã� P�8� ]Ë�U��M���E}�`�����Q�/  Y]Ã� P�8� ]���h�# d�5    �D$�l$�l$+�SVW� 1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�����������̋�U���S�]V�s35 W��E� �E�   �{���t�N�38�����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t����	  �E���|@G�E��؃��u΀}� t$����t�N�38�(����N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=� t h��H  ����t�UjR�����M�c	  �E9Xth W�Ӌ��f	  �E�M��H����t�N�38�����N�V�3:�����E��H����  �����9S�R���h W���	  ������U��V�uW3�;�u�����WWWWW�    ��������   �F����   �@��   �t�� �F��   ���F�  u	V�O  Y��F��v�vV����YP��M  ���F;���   �����   �F�uOV�����Y���t.V�����Y���t"V�������V�<��������Y��Y��H�@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�~���_^]�jTh� �����3��}��E�P�H� �E�����j@j ^V�  YY;��  ���5l��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@����   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j �(  YY��tV�M������l ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=l|���=l�e� ��~m�E����tV���tQ��tK�uQ�D� ��t<�u���������4���E� ���Fh�  �FP�%M  YY����   �F�E�C�E�9}�|�3ۋ���5�����t���t�N��r�F���uj�X�
��H������P�@� �����tC��t?W�D� ��t4�>%�   ��u�N@�	��u�Nh�  �FP�L  YY��t7�F�
�N@�����C���g����5l�<� 3��3�@Ëe��E�������������Ë�VW���>��t1��   �� t
�GP�L� ���@   ;�r��6������& Y�����|�_^Ë�U�����S3�V�u�E��]�]��]��F�> t��<at9<rt,<wt����SSSSS�    ������3��p  �E  ��M��]��E	  �M�3�AF�W:���  �Q� @  ;��.  ����S��   ��   �� �  ��tVHtG��t/��
t"����  9]���   �M�E�   ��   	U��   �E@��   �M@�   �E�   �   �E��   �E������E�E����E��   9]�uw�M �E�   �u��Tt\��tEHt1��t���  �E �  uF	}�L9]�u<�e������E�   �79]�u'	}��E�   �&�E �  u�M �  ��E   t3���M   F�:������9]���   �F�> t�jVhh� �8V  ������   ���F�> t��>=upF�> t�jhl� V�T  ����u���M   �Ajht� V�fT  ����u���M   �!jh�� V�FT  ����u���M   �F�> t�8t�����SSSSS�    �^������h�  �u�E��u�uP�Q  ����t3�� �E���M��H�M��X��X�X�H_^[��jh8� �n���3�3��}�j��'  Y�]�3��u�;5�,��   ����9t[� �@��uH� �  uA�F���w�FP�&  Y����   ���4�V�h���YY�����@�tPV����YYF둋��}��h��j8�  Y������9tIh�  � �� P�mH  YY����u�4����Y������� P�4� ���<�}�_;�t�g �  �_�_��_�O��E������   ������Ë}�j��%  Y���SVW�T$�D$�L$URPQQh�- d�5    � 3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C��T  �   �C��T  �d�    ��_^[ËL$�A   �   t3�D$�H3������U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�+T  3�3�3�3�3���U��SVWj j hS. Q�k�  _^[]�U�l$RQ�t$������]� ��U��V�uV�I���P��S  YY��t|������ ;�u3��������@;�u`3�@���F  uNSW�<���? �   u S�D  Y���u�Fj�F�X�F�F��?�~�>�^�^�N  3�_@[�3�^]Ë�U��} t'V�u�F   tV�����f�����f �& �f Y^]Ë�U��EV���F ��uc�z  �F�Hl��Hh�N�;t�$�Hpu��\  ��F;(t�F�$�Hpu�jU  �F�F�@pu�Hp�F�
���@�F��^]� �A@t�y t$�Ix��������QP��\  YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�����8*u�ϰ?�d����} �^[]Ë�U���x  � 3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������l�����u5�����    3�PPPPP������������ t
�������`p������
  �F@u^V����Y�H���t���t�ȃ�������������A$u����t���t�ȃ�����������@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw������ ��3��3�3������ j��Y������;���	  �$��; ��������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������\  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P��Z  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��������P�9X  Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������������/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V��  ������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�50��  Y�Ћ���������   t 9�����u������PS�5<�  Y��YY������gu;�u������PS�58�w  Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�[W  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u���������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�\U  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t�������B��������� Y���������������t������������������������� t
�������`p��������M�_^3�[������Ð�3 �1  2 ~2 �2 �2 3 I4 ��U���(  ���������5��=�f��f��f��f��f�%�f�-�����E ���E���E���������   ������	 ���   � ������� �������0� ��j�.  Yj �,� h�� �(� �=� uj�.  Yh	 ��$� P� � �Ë�U��V�5��5X� �օ�t!�����tP�5����Ѕ�t���  �'�� V�T� ��uV�  Y��th� P�� ��t�u�ЉE�E^]�j ����YË�U��V�5��5X� �օ�t!�����tP�5����Ѕ�t���  �'�� V�T� ��uV�   Y��th0� P�� ��t�u�ЉE�E^]��\� � ��V�5��X� ����u�5��e���Y��V�5��`� ��^á����tP�5��;���Y�Ѓ�������tP�d� ����  jhX� ������� V�T� ��uV�a  Y�E�u�F\�� 3�G�~��t$h� P�� �Ӊ��  h0� �u��Ӊ��  �~pƆ�   CƆK  C�Fh j��  Y�e� �vh�h� �E������>   j�  Y�}��E�Fl��u��Fl�vl��K  Y�E������   �b����3�G�uj�  Y�j�  YË�VW�� �5��������Ћ���uNh  j��  ��YY��t:V�5��5������Y�Ѕ�tj V�����YY�� �N���	V����Y3�W�l� _��^Ë�V��������uj�>  Y��^�jh�� �e����u����   �F$��tP�����Y�F,��tP����Y�F4��tP����Y�F<��tP����Y�F@��tP����Y�FD��tP�{���Y�FH��tP�m���Y�F\=�� tP�\���Yj�A  Y�e� �~h��tW�p� ��u�� tW�/���Y�E������W   j�  Y�E�   �~l��t#W��J  Y;=t��0t�? uW��H  Y�E������   V�����Y����� �uj��  YËuj��  YË�U��=��tK�} u'V�5��5X� �օ�t�5��5����ЉE^j �5��5�����Y���u�x��������t	j P�`� ]Ë�VW�� V�T� ��uV�R  Y�����^  �5� h`� W��hT� W����hH� W����h@� W���փ=� �5`� ��t�=� t�=� t��u$�X� ���d� ���= �5����\� �������   �5�P�օ���   �_  �5������5��������5��������5����u��������  ��teh�? �5������Y�У����tHh  j�   ��YY��t4V�5��5�����Y�Ѕ�tj V�y���YY�� �N��3�@��$���3�_^Ë�U��VW3��u��  ��Y��u'9�vV�t� ���  ;�v��������uʋ�_^]Ë�U��VW3�j �u�u��M  ������u'9�vV�t� ���  ;�v��������uË�_^]Ë�U��VW3��u�u��N  ��YY��u,9Et'9�vV�t� ���  ;�v��������u���_^]Ë�U��W��  W�t� �u�T� ���  ��`�  w��t�_]Ë�U���R  �u�hP  �5��D���h�   �Ѓ�]Ë�U��h|� �T� ��thl� P�� ��t�u��]Ë�U���u�����Y�u�x� �j�&  Y�j�C  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=d thd�E(  Y��t
�u�dY�@I  hP� h<� ����YY��uBh�K �`  �4� �$8� �c����=h Ythh��'  Y��tj jj �h3�]�jh�� �����j�B  Y�e� 3�C9��   ��E��} ��   �5\�����Y���}؅�tx�5X����Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5\�~������5X�q�����9}�u9E�t�}�}؉E����u܋}��h`� �T� �_���Yhh� �d� �O���Y�E������   �} u(�j�p  Y�u�����3�C�} tj�W  Y�����Ë�U��j j�u�������]�jj j ������Ë�V������V��
  V�6.  V�����V�R  V��Q  V��O  V�t  V��O  h�F ������$��^Ã=` u�B  V�5xW3���u����   <=tGV�:G  Y�t���u�jGW������YY�=���tˋ5xS�BV�	G  ��C�>=Yt1jS�����YY���tNVSP�tQ  ����t3�PPPPP�1��������> u��5x�����%x �' �T   3�Y[_^��5�������%� ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�xQ  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�P  Y��t��M�E�F��M��E���pP  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9`u�@  h  �VS��� ��,�5 ;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P������Y;�t)�U��E�P�WV�}�������E���H���5�3�����_^[�Ë�U�� ��SV�5�� W3�3�;�u.�֋�;�t�    �#�� ��xu
jX� �� ����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5�� SSS+�S��@PWSS�E��։E�;�t/P�9���Y�E�;�t!SS�u�P�u�WSS�օ�u�u������Y�]��]�W��� ���\��t;�u���� ��;��r���8t
@8u�@8u�+�@P�E��������Y;�uV�|� �E����u�VW�pN  ��V�|� ��_^[�Ë�V��� ��� W��;�s���t�Ѓ�;�r�_^Ë�V��� ��� W��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P��� �$��u]�3�@�P]Ã=PuWS3�98W�=� ~3V�5<��h �  j �v���� �6j �5$�׃�C;8|�^�5<j �5$��_[�5$��� �%$ �Ë�U��QQV����������F  �V\��W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ���=����;�}$k��~\�d9 �=���B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]Ë�U���� �e� �e� SW�N�@��  ��;�t��t	�У �`V�E�P��� �u�3u���� 3��� 3���� 3��E�P��� �E�3E�3�;�u�O�@����u������5 �։5 ^_[�Ë�U����M� � �	�` �H]� ��U��S�]V���� �C�F���CWt1��t'P�?  ��GW�,  YY�F��t�sWP�!J  ���	�f ��F_��^[]� �y �� t	�q�����YËA��u�� Ë�U��V��������EtV�u���Y��^]� ��Q�4� ��M  YË�U��V��������EtV�D���Y��^]� ��U��QSVW�5\�
����5X���}��������YY;���   ��+ߍC��rwW�N  ���CY;�sH�   ;�s���;�rP�u������YY��u�G;�r@P�u������YY��t1��P�4�����Y�\�u�������V�����Y�X�EY�3�_^[�Ë�Vjj �-�����V��������\�X��ujX^Ã& 3�^�jh�� ������-����e� �u�����Y�E��E������	   �E����������Ë�U���u���������YH]�jh�� �����e� �u;5@w"j��  Y�e� V��
  Y�E��E������	   �E������j��  YË�U��V�u�����   SW�=�� �=$ u�-E  j�{C  h�   �K���YY�P��u��t���3�@P���uV�S���Y��u��uF�����Vj �5$�׋؅�u.j^9t�u�G   Y��t�u�{���������0�����0_��[�V�    Y�����    3�^]Ë�U��E�(]Ë�U���5(����Y��t�u��Y��t3�@]�3�]Ë�U��� �EVWjY�8� �}��E��E_�E�^��t� t�E� @��E�P�u��u��u���� �� ��VW3��0�<��u����8h�  �0���"  YY��tF��$|�3�@_^Ã$�� 3����S�L� V��W�>��t�~tW��W�����& Y�����|ܾ�_���t	�~uP�Ӄ����|�^[Ë�U��E�4���8� ]�jh� �V���3�G�}�3�9$u�.C  j�|A  h�   �L���YY�u�4��9t���nj�����Y��;�u�	����    3��Qj
�Y   Y�]�9u,h�  W�!  YY��uW�M���Y������    �]���>�W�2���Y�E������	   �E�������j
�(���YË�U��EV�4���> uP�"���Y��uj�@���Y�6�4� ^]Ë�U��8�<k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ������   �L�5�� h @  ��H� �  SQ�֋L���   ���	P���@�L����    ���@�HC���H�yC u	�`����x�ueSj �p�֡��pj �5$�� �8��k��<+ȍL�Q�HQP��G  �E���8;�v�m�<�D�E���=L[_^�áHV�58W3�;�u4��k�P�5<W�5$��� ;�u3��x�H�58�<k�5<h�A  j�5$��� �F;�t�jh    h   W��� �F;�u�vW�5$�� 뛃N��>�~�8�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W��� ��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U����8�Mk�<������M���SI�� VW}�����M���������3���U��D����S�;#U�#��u
���];�r�;�u�<��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1�<�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t�D�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;�u�M�;Lu�%� �M���B_^[�Ë�U��EVW��|Y;lsQ���������<������<�u5�=�S�]u�� tHtHuSj��Sj��Sj���� ��3�[��<���� 	   �D����  ���_^]Ë�U��MS3�;�VW|[;lsS������<���������@t5�8�t0�=�u+�tItIuSj��Sj��Sj���� ���3������� 	   ��������_^[]Ë�U��E���u�����  ����� 	   ���]�V3�;�|";ls�ȃ����������@u$�a����0�G���VVVVV� 	   ������������ ^]�jh(� �����}����������4���E�   3�9^u6j
�S���Y�]�9^uh�  �FP�  YY��u�]��F�E������0   9]�t������������D8P�4� �E�������3ۋ}j
����YË�U��E�ȃ���������DP�8� ]�jhH� �W����M��3��}�j�����Y��u����b  j����Y�}��}؃�@�<  �4������   �u����   ;���   �Fu\�~ u9j
�K���Y3�C�]��~ uh�  �FP�  YY��u�]���F�e� �(   �}� u�^S�4� �FtS�8� ��@낋}؋u�j
����YÃ}� u��F��+4����������u�}��uyG�+���j@j �O���YY�E���ta�����l ���   ;�s�@ ���@
�` ��@�E������}�����σ�������DW�����Y��u�M���E������	   �E������j�R���YË�U���  �>C  � 3ŉE��EV3���4�����8�����0���9uu3���  ;�u'薾���0�|���VVVVV�    ����������  SW�}�����4�������ǊX$�����(�����'�����t��u0�M����u&�-���3��0����VVVVV�    虽�����C  �@ tjj j �u��@  ���u��  Y����  ��D���  �4����@l3�9H�������P��4�� ������ ���`  3�9� ���t���P  ��� ��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�m,  Y��t:��4���+�M3�@;���  j��@���SP�?  �������  C��D����jS��@���P�?  �������  3�PPj�M�Qj��@���QP�����C��D������ �����\  j ��<���PV�E�P��(���� �4��� ���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4��� ����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@����<  Yf;�@����h  ��8����� ��� t)jXP��@����d<  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4��� ���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4��� ���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  ��� ��;���   j ��,���P��+�P��5����P��(���� �4��� ��t�,���;����� ��@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0��� ��t��,�����@��� ��8������ ��@�����8��� ul��@��� t-j^9�@���u����� 	   �����0�?��@�������Y�1��(�����D@t��4����8u3��$�ķ���    �̷���  ������8���+�0���_[�M�3�^������jhp� 芹���E���u萷���  �u���� 	   ����   3�;�|;lr!�g����8�M���� 	   WWWWW�ն�����ɋ��������������L1��t�P�����Y�}���D0t�u�u�u�.������E������� 	   �����8�M���E������	   �E��
�����u�2���Y�jh�� 许���E���u衶��� 	   ����   3�;�|;lr耶��� 	   SSSSS�������Ћ����<����������L��t�P����Y�]���Dt1�u����YP��� ��u�� �E���]�9]�t�����M������ 	   �M���E������	   �E��)�����u�Q���YÃ%4 �����̋T$�L$��ti3��D$��u��   r�=0 t�:  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh�� �F���3ۉ]�j����Y�]�j_�}�;=�,}W�������9tD� �@�tP����Y���t�E��|(����� P�L� ���4�Q���Y���G��E������	   �E������j�<���Y�������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�� h�# d�    P��SVW� 1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����UV�uj�X�E�U�;�u�Q����  �6���� 	   ����  S3�;�|;5lr'�'��������SSSSS� 	   蕲��������Q  ����W�<�������ƊH��u������ǲ��� 	   �j�����wP�]�;��  ����  9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!�u�����[����    SSSSS�������4����M;�r�E�u�����Y�E�;�u�#����    �+����    ����h  jSS�u��4  ��D(�E���T,���AHtt�I��
tl9]tg��@�M�E�   �D
8]�tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4��� ���{  �M�;��p  ;M�g  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4��� ��u
�� ��uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�93  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@��� t��������u�ί��� *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u�_2  ���E�+]���P�uS�u�j h��  ��� �E���u4�� P�s���Y�M���E�;EtP让��Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E�É]�E�;���   �E�f����   f��tf�CC@@�E�   �M����;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4��� ��u
�� ��u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u��0  ��f�}�
tjXf�CC�E�9E�������t�@u��f� f�CC+]�]������� j^;�u�ǭ��� 	   �ϭ���0�i�����m�Y����]��\���3�_[^��jh�� 葯���E���u藭���  �|���� 	   ����   3�;�|;lr!�n����0�T���� 	   VVVVV�ܬ�����ɋ��������������L9��t�����;M�Au� ����0�����    �P�����Y�u���D8t�u�u�u�~������E���Ь��� 	   �ج���0�M���E������	   �E�������u����YË�U����h   �D���Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E��]�jh� �<����e� �u�u��� �E��/�E� � �E�3�=  �����Ëe�}�  �uj�l� �e� �E������E��.���Ë�U���0S3��E�VW���]��]��E�   �]�t	�]��E��
�E�   �]��E�P��4  Y��tSSSSS�������M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&�m�������P���j^SSSSS�0�٪�����   �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   t`;������E�   �E�E�   ��t����#M��x�E�   �@t�M�   �M�   �M��   t	}�� t�M�   ��E�   릨t�M�   ��������u������������    �   �E�=�� S�u��    �u�E�P�u��u��u�׉E���um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׉E���u4�6������������D0� ��� P�u���Y�I���� �t  �u��D� ;�uD�6������������D0� ��� ��V�2���Y�u��� ;�u�������    룃�u�M�@�	��u�M��u��6�+�����Ѓ������Y��Y�M����L��Ѓ���������D$� ��M��e�H�M���   �����  �Etqj���W�6�v0  ���E�;�u�p����8�   tM�6�P��������j�E�P�6�]����������u�}�u�E�RP�6�s.  ��;�t�SS�6�0  ��;�t��E���0  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   ��  �E�@�]���  �E��   �#�=   @��   =   �tw;���  �E�;��y  ��v��v0���f  �E�3�H�&  H�R  �E���  �E�   �  jSS�6��)  ���t�SSS�6��)  #���������j�E�P�6�w���������u�����tk����   �}�﻿ uY�E���   �E�;���   ���b������P���jSS�6�a)  ����C���SSS�6�L)  ��#����   �����E�%��  =��  u�6�F���Y�>���j^�0���d  =��  uSj�6�+.  �����������E��ASS�6�.  ����E�﻿ �E�   �E�+�P�D=�P�6�K��������������9}�ۋ������������D$�2M���0�������������D$�M�������
ʈ8]�u!�Et��ȃ���������D� �}��   ���#�;�u|�Etv�u��� S�u�E�jP�u������W�u��� ���u4�� P�5�����ȃ���������D� ��6�����Y�����6��������������_^[��jh0� 车��3��u�3��};���;�u襤��j_�8VVVVV�.��������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���j������E��E������   �E�;�t���v����3��}9u�t(9u�t�������������D� ��7�u���YË�U��j�u�u�u�u�u������]Ë�U���S�u�M�謱��3�9]u8]�t�E��`p�3���  �E�9Xu&�u�u�u��-  ��8]���  �M��ap��  9]u.�w���SSSSS�    �������8]�t�E��`p������  W�};�u.�A���SSSSS�    �ɢ����8]�t�E��`p������N  V�Mf�	�M�E�����D�M�ti9]u��D�]��  ��f����   �U�:�u�]��Z��f��f��E��f��M�f;prf;pwfp�6f;pr0f;pw*fp�$�U���Atf��  ����ʉM�f�u�f�����G�D�M�tH9]u�]��^��M:�t���f��f���G�M�f;Hrf;HwfH�6f;Hr0f;Hw*fH�$�U���Atf��  ����ʉM�f�M�f;�u!f;�t	9]�����8]�t�E��`p�3�^_[�����H8]�t��M��ap����U��j �u�u�u�������]Ë�U���S3�9]u3���   W�u�M��X����}�9_u&�u�u�u�Ó����8]���   �M��ap��   9]u+�=���SSSSS�    �Š����8]�t�E��`p������mV�u;�u+�
���SSSSS�    蒠����8]�t�E��`p������9�Ef� �M�E�����D8tA9]u�3��D8t_8]�t�E��`p�3�^_[�ËE� :�u3����f��f��E��f�����F�D:t 9]u3����M:�t�f����f�F��f;�uf;�t�9]�`�������H8]�t��M��ap�냋�U��j �u�u�u������]�U��SVWUj j h`� �u�^A  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�hh� d�5    � 3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �yh� u�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� ��Ë�U��E���u�˞��� 	   3�]�V3�;�|;lr譞��VVVVV� 	   �5�����3���ȃ���������D��@^]�-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�g���3��ȋ��~�~�~����~���� ���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  � 3ŉE�SW������P�v��� �   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R������C�C��u�j �v�������vPW������Pjj ��-  3�S�v������WPW������PW�vS�+  ��DS�v������WPW������Ph   �vS�+  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[蝓����jhP� �G���跺�����$�Gpt�l t�wh��uj ����Y���_����j�s���Y�e� �wh�u�;5(t6��tV�p� ��u�� tV�V���Y�(�Gh�5(�u�V�h� �E������   뎋u�j�8���YË�U���S3�S�M��~��������u��   ��� 8]�tE�M��ap��<���u��   ��� �ۃ��u�E��@��   ��8]�t�E��`p���[�Ë�U��� � 3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�0��   �E��0=�   r����  �p  ����  �d  ��P��� ���R  �E�PW��� ���3  h  �CVP�����3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�}����M��k�0�u���@�u��*�F��t(�>����E���,D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C��4Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95��X�������M�_^3�[蘐����jhp� �B����M��讷�����}�������_h�u�u����E;C�W  h   �Ǻ��Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�p� ��u�Fh= tP�2���Y�^hS�=h� ���Fp��   �$��   j�����Y�e� �C���C���C��3��E��}f�LCf�E�@��3��E�=  }�L�� 	@��3��E�=   }��  ��(
@���5(�p� ��u�(= tP�y���Y�(S���E������   �0j�m���Y��%���u �� tS�C���Y�ɗ���    ��e� �E������Ã=` uj��V���Y�`   3�Ë�U��SV�u���   3�W;�to=�th���   ;�t^9uZ���   ;�t9uP�ʑ�����   ��)  YY���   ;�t9uP詑�����   �)  YY���   葑�����   膑��YY���   ;�tD9u@���   -�   P�e������   ��   +�P�R������   +�P�D������   �9��������   �=(t9��   uP�o'  �7����YY�~P�E   ��(t�;�t9uP����Y9_�t�G;�t9uP�֐��Y���Mu�V�ǐ��Y_^[]Ë�U��SV�5h� W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�(t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5p� W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�(t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu��0tV�Y���Y��^�3��jh�� �ۖ���K�����$�Fpt"�~l t�4����pl��uj �y���Y�������j����Y�e� �Fl�=�i����E��E������   ��j�����Y�u�Ë�U��QV�uV�̐���E�FY��u�Q���� 	   �N ����/  �@t�6���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�<����� ;�t�0�����@;�u�u�����Y��uV�-���Y�F  W��   �F�>�H��N+�I;��N~WP�u�������E��M�� �F����y�M���t���t��������������H�@ tjSSQ�  #����t%�F�M��3�GW�EP�u�������E�9}�t	�N �����E%�   _[^�Ë�VW3����6訮����Y���(r�_^ËL$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v����j^SSSSS�0訑�������V�u�M������E�9X��   f�E��   f;�v6;�t;�vWSV�������̑��� *   ������ 8]�t�M��ap�_^[��;�t2;�w,衑��j"^SSSSS�0�*�����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p��� ;�t9]�^����M;�t����� ��z�D���;��g���;��_���WSV�1������O�����U��j �u�u�u�u�|�����]Ë�U����u�M�訞���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]��V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� jh�� �����M3�;�v.j�X3���;E�@u�Ώ���    WWWWW�V�����3���   �M��u;�u3�F3ۉ]���wi�=PuK������u�E;@w7j�����Y�}��u�����Y�E��E������_   �]�;�t�uWS�}�����;�uaVj�5$��� ��;�uL9=t3V萿��Y���r����E;��P����    �E���3��uj�{���Y�;�u�E;�t�    �������jh�� �͐���]��u�u�V���Y��  �u��uS����Y�  �=P��  3��}�����  j�����Y�}�S����Y�E�;���   ;5@wIVSP���������t�]��5V����Y�E�;�t'�C�H;�r��PS�u��  S�����E�SP�������9}�uH;�u3�F�u������uVW�5$��� �E�;�t �C�H;�r��PS�u��O  S�u��������E������.   �}� u1��uF������uVSj �5$��� ����u�]j����YË}����   9=t,V����Y��������e���9}�ul���� P����Y��_����   �@���9}�th�    �q��uFVSj �5$��� ����uV9t4V�{���Y��t���v�V�k���Y�����    3��,���������|�����u�ӌ������ P背���Y���ҋ�U��QQS�]VW3�3��}�;�@t	G�}���r���w  j�H%  Y���4  j�7%  Y��u�=��  ���   �A  h�� �  S��W��  ����tVVVVV袊����h  ��Vj �� �� ��u&h�� h�  V�  ����t3�PPPPP�^�����V�����@Y��<v8V�������;�j��h�� +�QP�  ����t3�VVVVV�������3�h�� SW��  ����tVVVVV��������E��4�DSW�  ����tVVVVV�҉����h  h�� W�"  ���2j��@� ��;�t$���tj �E�P�4�D�6�7���YP�6S��� _^[��j��#  Y��tj�#  Y��u�=�uh�   �)���h�   ����YY�jh�� �Ό���>����@x��t�e� ���3�@Ëe��E������#  �����h�� �E���Y��Ë�U��E��������]Ë�U��E��V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5��Y���Y�j h� �"���3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�������}؅�u����a  �����`�w\���]���������Z�Ã�t<��t+Ht貉���    3�PPPPP�8�����뮾���������
�����E�   P蕥���E�Y3��}���   9E�uj舮��9E�tP覻��Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.���M܋����9M�}�M�k��W\�D�E����������E������   ��u�wdS�U�Y��]�}؃}� tj �4���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��Ċ��Ë�U��E��]Ë�U��E�]Ë�U��MS3�VW;�t�};�w�C���j^�0SSSSS�̇�������0�u;�u��ڋъ�BF:�tOu�;�u�����j"Y�����3�_^[]Ë�U����u�M��ȕ���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]��U��WV�u�M�}�����;�v;���  ��   r�=0 tWV����;�^_u^_]��!  ��   u������r*��$�D� ��Ǻ   ��r����$�X� �$�T� ��$�ؚ �h� �� �� #ъ��F�G�F���G������r���$�D� �I #ъ��F���G������r���$�D� �#ъ���������r���$�D� �I ;� (�  � � � �  � �� �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�D� ��T� \� h� |� �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��� �����$��� �I �Ǻ   ��r��+��$�� �$��� ��� � @� �F#шG��������r�����$��� �I �F#шG�F���G������r�����$��� ��F#шG�F�G�F���G�������V�������$��� �I �� �� �� �� �� �� Ĝ ל �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��� ��� �� � � �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��jh0� ����j�u���Y�e� �u�N��t/���E��t9u,�H�JP�X~��Y�v�O~��Y�f �E������
   �
���Ë���j�@���Y�����������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����jhP� ����3��]3�;���;�u�����    WWWWW苂��������S�=Pu8j�<���Y�}�S�e���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5$��� �����؄���3��]�u�j�
���Y������U��WV�u�M�}�����;�v;���  ��   r�=0 tWV����;�^_u^_]��  ��   u������r*��$�T� ��Ǻ   ��r����$�h� �$�d� ��$�� �x� �� ȟ #ъ��F�G�F���G������r���$�T� �I #ъ��F���G������r���$�T� �#ъ���������r���$�T� �I K� 8� 0� (�  � � � � �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�T� ��d� l� x� �� �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�� �����$��� �I �Ǻ   ��r��+��$��� �$�� �� (� P� �F#шG��������r�����$�� �I �F#шG�F���G������r�����$�� ��F#шG�F�G�F���G�������V�������$�� �I �� �� �� �� ġ ̡ ԡ � �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�� �� � � � ,� �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U���� 3ŉE�V3�95tO�=8�u�x  �8���u���  �pV�M�Qj�MQP� � ��ug�=u��� ��xuω5VVj�E�Pj�EPV��� P��� �8���t�V�U�RP�E�PQ��� ��t�f�E�M�3�^�u�����   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M�������E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p��� ���E�u�M;��   r 8^t���   8]��e����M��ap��Y����|}��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p��� ���:���뺋�U��j �u�u�u�������]Ë�U��QQ�EV�u�E��EWV�E��b������Y;�u��|��� 	   �ǋ��J�u�M�Q�u�P�� �E�;�u�� ��t	P��|��Y�ϋ�����������D0� ��E��U�_^��jhp� �~������u܉u��E���u�|���  �r|��� 	   �Ƌ���   3�;�|;lr!�c|���8�I|��� 	   WWWWW��{�����ȋ��������������L1��u&�"|���8�|��� 	   WWWWW�{����������[P辺��Y�}���D0t�u�u�u�u�������E܉U���{��� 	   ��{���8�M���M���E������   �E܋U���}����u�����Y��������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh�� �_|���e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E��a|��Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[�������03�Ë�U���SVW3�jSS�u�]��]��l����E�#��U���tYjSS�u�P�����#ʃ����tA�u�}+����   ;���   �   Sj�� P��� �E���u�*y���    �y��� _^[��h �  �u�  YY�E���|
;�r�����P�u��u�!��������t6�+��xӅ�wϋu��u��u�F  YY�u�j �� P�� 3��   �x���8u�x���    ����u��;�q|;�skS�u�u�u�U���#�����D����u迶��YP�� �����H��E�#U���u)�>x���    �Fx������ ��u�#u��������S�u��u��u�����#���������3��������U��V�uV�F���Y���u��w��� 	   ����MW�uj �uP�� �����u�� �3���tP��w��Y����������������D0� ���_^]Ë�U��S�]V�u�������������0�A$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��EV3�;�u�v��VVVVV�    �9v����jX�
�t�3�^]Ë�U���S3�VW9]��   �u�M��N���9]u.�av��SSSSS�    ��u����8]�t�E��`p������   �};�t˾���9uv(�"v��SSSSS�    �u����8]�t�E��`p����`�E�9Xu�uW�u��  ��8]�tD�M��ap��;�E� �M�QP�  �E����M�QP�  ��G�Mt;�t;�t�+����3�_^[�Ë�U��V3�95�u99uu�u��VVVVV�    �u���������'9ut܁}���w�^]�E  V�u�u�u������^]Ë�U��E��t���8��  uP�o��Y]Ë�U���� 3ŉE�SV3�W��9u8SS3�GWh�� h   S�� ��t�=��� ��xu
�   9]~"�M�EI8t@;�u�����E+�H;E}@�E�����  ;���  ����  �]�9] u��@�E �5�� 3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�v  ��;�t� ��  �P覣��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5� SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�  ��;�tj���  ���P����Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�� ��t"SS9]uSS��u�u�u�VS�u ��� �E�V����Y�u������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�  Y�E���u3��!  ;E ��   SS�MQ�uP�u �-  ���E�;�tԋ5� SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�  ��;�t����  ���P�Ρ��Y;�t	� ��  �����3�;�t��u�SW�H������u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��|  ���u������#u�W����Y��u�u�u�u�u�u�� ��9]�t	�u��l��Y�E�;�t9EtP� l��Y�ƍe�_^[�M�3���h���Ë�U����u�M��G���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ� 3ŉE��SV3�W��;�u:�E�P3�FVh�� V�� ��t�5�4�� ��xu
jX�������   ;���   ����   �]�9]u��@�E�5�� 3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�  ��;�t� ��  �P����Y;�t	� ��  ���؅�ti�?Pj S�f�����WS�u�uj�u�օ�t�uPS�u�� �E�S������E�Y�u3�9]u��@�E9]u��@�E�u�0  Y���u3��G;EtSS�MQ�uP�u�X  ����;�t܉u�u�u�u�u�u�� ��;�tV�j��Y�Ǎe�_^[�M�3���f���Ë�U����u�M��H}���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v�i���v�i���v�i���v�yi���v�qi���v�ii���6�bi���v �Zi���v$�Ri���v(�Ji���v,�Bi���v0�:i���v4�2i���v�*i���v8�"i���v<�i����@�v@�i���vD�i���vH��h���vL��h���vP��h���vT��h���vX��h���v\��h���v`��h���vd��h���vh�h���vl�h���vp�h���vt�h���vx�h���v|�h����@���   �h�����   �~h�����   �sh�����   �hh�����   �]h�����   �Rh�����   �Gh�����   �<h�����   �1h�����   �&h�����   �h����,^]Ë�U��V�u��t5�;�tP��g��Y�F;�tP��g��Y�v;5�tV��g��Y^]Ë�U��V�u��t~�F;�tP�g��Y�F;�tP�g��Y�F;�tP�g��Y�F; tP�|g��Y�F;tP�jg��Y�F ;tP�Xg��Y�v$;5tV�Fg��Y^]Ë�U��ES3�VW;�t�};�w�l��j^�0SSSSS�:l�������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��jl��j"Y����3�_^[]���������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w��k��j^�0SSSSS�]k��������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����Zk��j"Y���������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^��j�͍��YË�U���VW�u�M���x���E�u3�;�t�0;�u,��j��WWWWW�    �_j�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�
  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&�6i���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9�uh�P������]Ë�U���SVW蹄���e� �=$ ����   h�� ��� �����*  �5� h�� W�օ��  P�����$|� W�$��P�����$h� W�(��P�ك���$L� W�,��P�ă��Y�4��th4� W��P謃��Y�0�0;�tO94tGP�
����54�������YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9�(;�t0P躃��Y��t%�ЉE���t�,;�tP蝃��Y��t�u��ЉE��5$腃��Y��t�u�u�u�u����3�_^[�Ë�U��MV3�;�|��~��u���(������g��VVVVV�    �f�������^]Ë�U���(  � 3ŉE��0Vtj
����Y������tj����Y�0��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�Z�������������(�����0���j ǅ����  @��������,����,� ��(���P�(� j�����U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]�3�PPjPjh   @h�� ��� �8á8V�5� ���t���tP�֡4���t���tP��^Ë�U���SV�u�M���q���]�   ;�sT�M胹�   ~�E�PjS�  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P����YY��t�Ej�E��]��E� Y��qc��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�������$���o������E�t	�M�����}� t�M��ap�^[���������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���� 3ŉE�j�E�Ph  �u�E� � � ��u����
�E�P��  Y�M�3��Y���Ë�U���4� 3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5�� �M�QP�֋�� ��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��������YF;�~[�����wS�D6=   w/�  ��;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�#���Y;�t	� ��  ���E���}�9}�t؍6PW�u�藫����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u��� ��t`�]��[��� 9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�����YY�E�;�t+WWVPV�u�W�u��;�u�u��Q[��Y�}���}��t�MЉ�u�����Y�E��e�_^[�M�3���W������Q�L$+ȃ����Y����Q�L$+ȃ����Y������U��j
j �u������]Ë�U���S�u�M��9n���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�I���YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�h����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%P� ��`� ������                                                                                                                                                                                                                                                                                                        �  .�  D�  ��  ��  ��  ��  ��  ��  ��  
�  &�  D�  X�  p�  ��  ��  ��  ��  ��  ��  ��  �  �  �  *�  4�  L�  \�  t�  |�  ��  ��  ��  ��  ��  �  �  "�  0�  J�  Z�  p�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  .�  :�  b�  p�  |�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  *�  :�  J�  \�  n�      d�  r�                  �! !P �� ��         � \"                     ��R       f   P�  P�  bad allocation  Can't load anima dlls   .cdl    Anima.C4D12 \   found programPath %s
   PATH    Anima.xml File not found!
  Anima.xml File not found!   an(i)ma StartupError    r   Anima.xml   c4d_main        �� ' O ccs UTF-8   UTF-16LE    UNICODE ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          � EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       8� O O Unknown exception   L� FO csm�               �        	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL   Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        0� (� � � � �� �� �� �� �� �� � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� |� x� t� p� l� h� d� `� \� X� T� P� L� H� D� @� <� 8� 4� 0� ,� (� $�  � � � � �� �� �� �� �� �� x� X� 8� � �� �� �� �� l� P� @� <� 4� $�  � �� �� �� �� �� x� P� (� �� �� �� �� l� @� $� �� CONOUT$ SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    H                                                            ��    RSDS��K,'22N�S�PbXn   C:\Lavoro\anima\sdk\src\Anima.Plugin\C4D\obj\AnimaWrapper12_Win32_Release.pdb                ��            �� �� �             ����    @   �� 8         ����    @    �            0� �                 8  �             �`�            p� x�     �        ����    @   `�             �#  �-  h�                      ����    ����    ����    �     ����    ����    ����    �     ����    ����    ����    �     ����    ����    ����    J     ����    ����    ����� �          l�    x� ��          ����       N     8     ����       �N ����    ����    ����    &     ����    ����    ����    �     ����    ����    ����    �         w ����    ����    �����( �(     ����    ����    ����    -     ����    ����    ����    @? ����    O? ����    ����    ����    A ����    A ����    ����    ����    |F     ����    ����    ����    �P     ����    ����    ����    �P     ����    ����    ����    �S     ����    ����    ����    �`     ����    ����    ����    �b         �a ����    ����    ����    �j     ����    ����    ����    yk     ����    ����    ����    �l     ����    ����    �����m �m     ����    ����    ����    �t     ����    ����    ����5u Lu     ����    ����    ����    ,}     ����    ����    ����    ��     ����    ����    ����    o�     ����    ����    ����    ߌ     ����    ����    ����    \�     ����    ����    ����    ��     ����    ����    ������ ��     ����    ����    ����    ��     ����    ����    ����    ��     ����    ����    ����    ʞ     ����    ����    ����    ϥ     ����    ����    ����� *� ��          V�   �  �          ��  (�                      �  .�  D�  ��  ��  ��  ��  ��  ��  ��  
�  &�  D�  X�  p�  ��  ��  ��  ��  ��  ��  ��  �  �  �  *�  4�  L�  \�  t�  |�  ��  ��  ��  ��  ��  �  �  "�  0�  J�  Z�  p�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  .�  :�  b�  p�  |�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  *�  :�  J�  \�  n�      d�  r�      �LoadLibraryExA  �GetModuleFileNameA   GetProcAddress  KERNEL32.dll  �MessageBoxA � GetActiveWindow USER32.dll  �GetCurrentThreadId  oGetCommandLineA �GetLastError  �HeapFree  C CloseHandle -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent � EnterCriticalSection  �LeaveCriticalSection  �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA � DeleteCriticalSection �RtlUnwind �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �InterlockedIncrement  �SetLastError  �InterlockedDecrement  !Sleep ExitProcess JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW zWideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapAlloc ZRaiseException  TVirtualAlloc  �HeapReAlloc �SetStdHandle  �WriteFile �GetConsoleCP  �GetConsoleMode  AFlushFileBuffers  MultiByteToWideChar hReadFile  �InitializeCriticalSectionAndSpinCount x CreateFileA [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �LoadLibraryA  �HeapSize  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW �SetFilePointer  �SetEndOfFile  #GetProcessHeap  �LCMapStringA  �LCMapStringW  =GetStringTypeA  @GetStringTypeW  �GetLocaleInfoA      ��R    ��           ��  ��  ��  p  ��    AnimaWrapper12.cdl c4d_main                                                   �� ��         N�@���D�� 4�     .?AVbad_alloc@std@@ 4�     .?AVexception@std@@                                      	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����
                                                          �� �� ���������F          x   
   �� �� 4�     .?AVtype_info@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                      �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    � ����C                                                                                              (            (            (            (            (                              �         � �� � (0   0 P� P� P� P� P� P� P� P� P� P�    h�    <� 	   � 
   x�    L�    �    ��    ��    ��    l�    4�    ��    ��    ��    P�     � !    � "   �� x   p� y   `� z   P� �   L� �   <�         ��                             � � 0� ,� (� $�  � � � � �  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� x� p� h� \� T� H� <� 8� 4� (� � � 	         (.   �         �   .                 ��������    �p     ����    PST                                                             PDT                                                             P�����        ����        ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                                                                                                                                                                                                                                                                                                                                                                                                                                             �   00:0E0b0o0�0�0�0�0�0�0�011K1�1�1�1�1�1�1 222%2+20282B2y2~2�2G3�455;5B5�5N6�6^7i7�8�8�8�8.9F9N9T9�9�9�9�9::r:�:;;;1;`;�;�;�;�;�;�;�;4<:<K<u<�<�<�<�<1=`=�> ??.?}?�?�?      �   �0�0�0�0�0�0'1C1f1y1�1�1�1�1�1�1�122 2-2Q2c2q2�2�2�2�2�23%3T3]3z3�3�4�4�4�4;56!6z6�6�6�6�6>7F7�7�7�7�78B8T8�8�8�8�89"9�:;:;Z;�;�;<<H<X<�<�<�<�<�<�<1===I>�>�>i?q?�?�?   0  �   x0181^1�1�1�175'6�7�78�9�;�;�;�;�;�;�; <<<<"<(<.<5<<<C<J<Q<X<_<g<o<w<�<�<�<�<�<�<�<�<�<�<�<�<�<�<===#=/=D=K=_=f=�=�=�=�=�=�=�=�=�=>>>&>,>5>A>O>U>a>g>t>~>�>�>�>�>�>�>�>?^?d?�?�?�?�?�?   @  T  h0�0�0�0�0!11171C1I1Y1_1t1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122222!2'2,22272F2\2g2l2w2|2�2�2�2�2�2�2�2�2�2/383D3{3�3�3�3�3�34484S4Y4b4i4�4�4�4555%5/565A5J5`5k5�5�5�5�5�5�5656:6E6J6h6�67	77P7Z7�7�7�7�7�7�9�9�9�9�9�9$:*:@:K:b:n:{:�:�:;;M;f;u;z;�;�;�;�;�;�;�;<<<(<4<=<E<O<U<[<}<�<�<==�=>>'>/>7>C>g>o>�>�>�>?;?r?}?�?   P  �   090>0U0�0�0
1101g1x1�1�1292H2O2Y2�2�2�2�2�2�2�2�2�2343�3�3�3�3?6M6S6m6r6�6�6�6�6�6�6�6�6�6�6�6	7777'7-777>7R7Y7_7m7t7y7�7�7�7�7�7�7�7<8�;�;<=<w<�<�>�>�>�>�>�>?H?X?s?�?�?�? `  x   50Q0�0�0�0�0�0<1N1�1�1�122]2�23�3�3�4�4N5�6�7�8�8�89,9�9�9,:�:�:�:0;:;�;�;<.<:<a<n<s<�<H=M=_=}=�=�==>s>�?   p  T   �0�0r1�1�12�2�2�3�3�3%4�455,5\57�7�78818D8V8�8�8�;�;�;<8<C<Z<<�<K=   �  �   T1�1�1=2W2`2�2�2E3�3�355W5d5n5|5�5�5�5�5�5�5�5626i6�6�6!7>7�7�78�8�8�8�8�8�8�8�89.979=9F9K9Z9�9�9�9�9�:�:;d;�;�;a<x<�<�<�=�=W> �    0:0h1�1�12%212�2�2�2\3b3�3�3�3 444:4F4�4�4�45535<5C5L5�5�5�5�566.6@6d6�6�6�6�6�6�6�6�6#717x7}7�7�7�7�7�7�7N8W8]8�8�8�9/:H:O:W:\:`:d:�:�:�:�:�:�:�:�:�:�:�:>;D;H;L;P;�;�;�;�;�;�;�;<;<m<t<x<|<�<�<�<�<�<�<�<�<�<�<8=X=]=;>s>�>�>
???X?_?g?l?p?t?�?�?�?�?�?�?�?�?�? �  �    00N0T0X0\0`0�0�0�0�0�0�0 1!1K1}1�1�1�1�1�1�1�1�1�1�1�1�1�1N2\2d2q2�2�2�2�2�2�2�2�2 3�344�4�4�4505�6�78"8�8�8 9-9�9�9�9�9�:�;I<[<h<t<~<�<�<�<�<�=8>[>�>�?   �  �   20<0T0[0e0m0z0�0�0J1�1�3�3�34$464H4Z4l4~4�8�8�8�8�8�8�8
999%949:9H9Q9`9e9o9}9�9�9�96:=:C:s:~:�:e;r;�<�<===!=�>�>?<?I? �     (070�2�2�2�2 �  (   @1D1H1L1X1\1\2`2d2�2 34440444 �  (  @:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;D<H<�<�<�<�<�<�< ===,=0=D=H=X=\=l=p=x=�=�=�=>8>T>X>`>h>p>t>|>�>�>�>�>�>??,?0?P?p?|?�?�?�?�? �  @    0 0@0`0l0�0�0�0�0�01$1(1H1h1�1�1�1�122(2H2h2�2�2�2     �    000080�1�1�4�4�4�4�4�4(; <�<�<�<�<�<�<�<�< ======= =$=(=,=0=4=8=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= > >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ?????�?�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              