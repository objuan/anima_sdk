MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       d��= �n �n �n�� n!�n;&n8�n;n��n)�+n%�n �n|�n;nd�n;#n!�n;%n!�nRich �n        PE  L ���R        � !
  �  �     ��                             �    �9
  @                   �� [    <      �                   0 �B  @~                                            L                           .textbss�                        �  �.text   ��  �  �                   `.rdata  B  p  D  �             @  @.data   I   �     �             @  �.idata  �        	             @  �.rsrc   �         	             @  @.reloc  �M   0  N   	             @  B                                                                                                                                                                                                                                                                                ������ �a �� 闲 ��h �Gf �� �C� �.� �9� �s �� �Z �5� �`�  ��, 鶲 ��k �7 釟  �¡ �}� �� �#U �.8 �)L �d[ �� 銵 �5- �$f �K\ 馄  �;g �z 鷮  �r� �ͭ ���  飰 鮄 �� ��@ ��� �ښ �r 鐁 ��  �VC �Q �l� �p  �Ҕ �̈́ �n ��b �^�  �#� ��� ���  �r �I ��W �ۮ �vt �1B �`  �� �h  ��  �8�  �C�  �~h �� �d� �_W  �z` ���  �Ѓ �{� ��  顆  ��  ��! �a � �h�  郬 �= ��y �d7 ��d �� �%� � � �۱  �{ � �H �� �R\  �� ��( �& �	 �f ��� �?� �
> ���  �p�  �;( �� �f  � �A ��! �=_ ��p �S �� ���  �d �o ��? �� � �  ���  �v� �1u �y �N �b� �n �XB ��h �. �YA �$ 鯗 �گ �5�  �Zd �K�  閑 �Az �zc �z �T �]� �x� �� �>�  �i� �t� �O�  �ʪ  �E9 �� �� ��P �b �5 �7O ��� ��� �Q  �s  �v �)d  �( ��i �c �� � �  �;y ���  �Q% �= ���  �b{ �M�  �H, �s= �~� �YJ �z �x ��D �O �`�  �k� �~ ��c ��v � �,b �� �Z �S� �ι  ��  ��@ �n �Zq 鵥  �Д  鋳 �O ��G 鬝 �G> �3 �}� �Pb �Ӝ �>� �b ���  �Ϥ  ��=  �� �М ��a �6 ��l  �? �7j �r� 鯅 �= �C� �x  �9L �D �Ol  �:� �%� 鰔 �+R ��  ��B �,; 闲  ��b �=� ��  �S� ��E �O �, �?� �J�  ��  �P� �[` �v� �� ��u �w1 ���  �]A �H� �� �a �	O �ī 鯩 ��{ �U� ��M  �( ��� �1F �\�  ��w �BQ ��p  �: �c� �! �		 �4�  �O@ �z< ��� ��� ��i �} �F �\ �ws �B= ��\ �za �y ��r �P �t �" �3 �5r ��O 鋨  �[ �6 ��  闟 ��[ ���  �د  �CU �< �y\ �] ��  �
� � ���  ��s �� �� �� �� �4 �-�  �(� �Ӎ �>X �98 �$c  ��� �_ ��O ��6 �a ��� �ac �\z �7r �� ��G �xN �3�  �
a �� ��� �L  �* ��) 鰃 ��c �V� ��  �,a �] � ��� �,_ �] �.I �Y �X �- �` �, ��� ��u  ���  �A� �M �s 颩 魧 �Xy  � �` �ٲ  ��� 韈 �
� �c` 逤  �ˏ �� �A� �l�  �'t  � �` �� �> 龐 �	 �D�  �3_ �� �e� � ��� �V_ �ч �\� ��  �R� �M� 鈼  ��� �ޚ �i �� �_ �4 �E
 ��x �k�  �6�  �!� �w �g� �b� ��H ���  �c2 �6 �)�  ��1 �K^ �� �5� �i� �� �& �Q�  �T  �� ��$ �� �h$ ��| �� �9�  ��t 鯤  �JZ �}� �P1 ��� � �� ���  �G� ��^ �ݵ �H� �6 �< �i�  �� �/9  ��: �U� � �+�  �� �q� � ��  �Ҳ  �}�  ��� ��� �` �Y� � �F ��X ��� � �[ �V�  �G �~Z � �"z �]t � �c �� �9� �$  ��7 ���  ��f �� �+e �v� �� ��  �� �bA ��  �H} �c� �� �i�  ��s �< �i �Յ � �\ ��U �Q �l� �7A �P ��[ �s  ��h  �b\ ��t �T� �� ��� ��8 ��< �+� 醭 鑑 �̛ �'] ��d �]x �h7  ��  �.� �� ��� �7  �JD ��= �w �E  �E �? �l� �wm �� ��  �H' ��( �.Z �)m �tV �?�  �@ �5�  �� �;:  ��� ��m �[ �7i �r? ��� �[ ��- ��0 ��P �L  �/M  � ��  � 4 ��@ �F� ��| �D �7 �� �]| �; �  �Μ  �y �J �O`  �ZN  �� �P� 雉 �&� �� ��  ��  �z ��  �h�  �c� �.n �9 �T� �� �� ��� �PN �S �Vp �1% �|�  �W<  �"K �& ��z �� �. �IT �4�  �? �*�  �e, �[ �K �V� �� ��Z �� 邤 ��b ��  �Z 龧  ��c �T� � �
� �� ���  ��  ��Y �Q0 ��  �| �H �=T ��  �v �� �9 � �v �f �I  �9 點 ��  ��  �XZ �'! �H �CZ �(C  �R �>' �)�  �6 �*W �ʖ �Z 鰄 �kc ��w �A4 �<P  �� ��  � �� �C� �P �Y 鴜 ��� �:I ���  ���  �k7 �F� �5Z �,K �'  ��g �� ��/ 飹 �� �y ��  �_Y  �:�  �, ��  ��r �v� �Q( ��P �U ��� ��  ��  �l ��  ��� 锢 �_r �Z� �U� �pG 髾  ��E �!�  �<  �'W  � �-� �h� �#� �.e �u �R �+ �J ��k ��  �kP  � �� �,� �� �X �- ��  ��i �.� �> �T4 ���  �JP �u. �  �+� �� �!�  ���  �g]  �r4 ���  ��U �m �>I � �r 鿋 �z� �UD �`� ��7 ��� �W �K �R �b�  �-� �h 鳔 �G  ��K �1 �1X �Zo ��}  �G  � �6� �� �� ���  钁 ��  ��f �4 �.a ��H �� ��� �zp  �H �0� 黩  �F� �S ��0 駱  �� ��g �{ �#�  �w  �d  ��� ��5  �z5  �� �`F �y �F� ��� �|= ��  ��  魬 �� �ӻ � �ih 鴾 �o/ �*i �~ ��m ��: �� ��� �̵  �gr  �~� 魤  ���  �S�  ��> �B �x ��  �
j  �C �`7 �J �&� �) �|� �'� �r�  �� 鸟 �#�  �^~ �I\  锢 �� �� �5u �@� ��V �s �qF  鬟 �GP �c ��U �ȓ �3$ �x �f �
 �O2 ��� �E�  �Z  �/ � �A�  �l5 �� 鲒 ���  阛 铑  �M �yf �` ���  �Zl �e ��  �V �ֿ  ��  ��j �� �� �L ��  ���  �U ��� �t�  �[T �Zs �%�  ��� 髜 �F8 �q�  �d  ��  �r} ��s �X5 �cb �^a �y� �t� ��  �z�  �5` �n �[ ��T �A� �0 � ��  �- �h� 鳓 �.j �i~ �$�  �_� �J� �V �� ��S �f�  ��v �|� �' �B? �A �� 飢 �^r �n �Đ  �qS �ʸ ��S �0 ��� �f& ���  �LI  �h 還 �y  �a  ��} �.� �	} �- ��  �ZT ��p �x ��>  �� �!�  �o  ��( �RR �ɿ � �s" �n� ��  �D�  ��S �J� � �`�  �Y �Fp �qE �l_ ��c ��  �]�  �Xb ��0 �>� ��{ �` ��  ��d �5m �`�  �{: ��X �q�  �G  �7� �B �T  �؊ �� �~q � ��� �ߒ  �
g � �P� �� �6P ��\ ��  �} �Bk ��b ��: ��R �.k  �9.  �� �?� �J# ��� �8 ��� �&� �� ��M �" �Bd �}K  ��] �c�  �`R �� �� �[ �Ze �U< ��G �k�  �Ơ  �% �V �l ��a ���  �R �Q �> ��� �4A �
 麃 �" �9 �[� �> �F  ��N �T �r7 靹  �N �3 �N �N ��P �n �Ji ��� � ; ��  ��;  �Q �� �'�  � �]� �x�  �c� �� �f �� �' �z� �$ �`? �+� �f�  鱴  �<> �7 �b� ��  ��H �sK �^� ��  �4�  �O�  �w �� � �� �6] �a�  �7  �Wc �R� ��0 �(B �C ��c  �I?  � 騎 �Z� ��  �U �K � ��� �G �'P  ��� �$ �k �cx ��� �Y� �Ԛ �o/ �j�  ��  ��� �I �O �!� ��� �1 ��  ��� �=  郜 �^l �I�  �$�  �" ��`  �e4  ���  �P �r �o ��9 �7�  �r �^ �h@ �c �.u  �Y� �4� �" ��} �e ��s  �[K  �] ��� �n ��t �"f �}h �" �Y �i ��4  �W �/�  �*K �U ���  �ۊ �} �Q�  �</  �C  �� ��9  �(! ��� �^] �)� ��j �+O �- �%F  這  �KH ��K �A! �l� �C � 齽  �x� �z �! �N ��� �� ��J �u �[  �[G  �VN �1 �s �g5 ��q �]� ��N �s�  �+ 驁 �� �K �h ��N ��e  ��  �65 �!� ��  �M �b? �* �(� 飈  ���  �I2  �hM �9  �
� �� �@L �;P  �v� �A� �\� 闵 �� �}� �; �1 �W ��� �� �o�  �j� �U� �pH  �k& �Fz �Q� �,� �g�  �r} �]� �e �� �s ��| ���  �o �A  �O ��> �{�  �6M ��� �<� � �bX ��� �83 �S  �~ �i�  ��d �?� ��& ��e �@] �;f � �qz � �W: � �}P 鸹 �s� �v  �y, �� ��6 ��g �E ��' 鋒 ��L �q�  ��  �L �a �=Q �xe �#�  ��  ��< �$� �J � �eQ �� �L ��w  ��a  �<� 闩 �r( �i  �VL �* ��L �� �$\ �_ �Z �P �`� ��; ��  �� �,t �Gg �a ��) �w �#� �a �IE �L �u  ��a ��  �zL �?L �\  �Au �̶ �� �Y ��,  �H� �# �>� �)p  �4�  ��&  �� �u� �TL �* ��  ��V  � � ��+  ���  �(�  �C� �^8  �K ��k �O]  �} �Ue ��� �� ��  ��| ���  �� �F �H � ��  �>� �i$ �$� �W �*� �Ş �I �k�  �v� ��& �LF 駧 �B� ��^ ��  ��H  �K ��� � 鿝  �J � ��� �۳  �� ��l 鬶 �� �2  齦 �h �S+  ��)  �U 鄩 ��' �6 ��I �`5 ��  �$ �� �� �� ��a �x  �Hz ��  �N� ��b �m  ��c �j� �- �0�  �ۉ �v� �'� �$ ��� �R� �=� �6J �3� �.�  ��q  �F  ��7 ��R �+ �6I �[C �6 �!� �l/  ��H �bw �v  �� �S� �^�  �)F  ��  �  隒  �� �@I ��7 ��+ ��V �B �g� �� �� �k  �C�  �N� ��  �TL  �uH ��� �u6 �8 ��� �� ��  �<I ��y �2� �Ma  �Ht ���  �~�  ��y �� �? ��  �I 鐊 �{� �vW  ��V  ��B  駅 �� ��  阔  � �� �ك �4L  �/� 銎 � �@ �+} �6& ��� 錗 �7� �D ���  �@ ��_ �n� �y�  �t� �Op �ʁ �U� �0 �+� �k �q �' �G  �2� � �� �C� �N� �	C �Ԙ �; �y �E� �`� �;w  �# �q� ��� �W� �R� ��H �H�  �yH �.[ ��� �v �n  ��^ �5f ��w �+Z �� � ��F �w� �H �-" �xK  �. 鮬 鉎 �@ �_�  �ZD  �B �p� �;� �� ��z  �|� �'" �� �]; �8� �Sw  ��q �Y  ��G ��; ��  �5^ �� � �i �у �M  �7� �"� �� � �c; �~�  ��V �dY �a  �*D  �%X �C �� ��  ��W  錻  �<  �"� �� �� �sp  ��T ��� �6 �� ��  �� ��@ 髢 ��W ��8  � �Gt �2�  �]� �F �\ �� �9� ��y �O� �E 饂 ���  �o � �?  �\� �w/ ��f  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��]�S����������U��Ejj j P�������]����������U��Ejj j P�������]����������U��]������������U��EHu�E�M�����   ]� �������������U����  ���3ŉE��=� �  VWjj j h  �R��������h  VP�Pj\V�{�����+��OQ������VR�l�����������Ƅ=���� H�H@��u��T��X��f�\��P������Rf�H�{���V����������hP�P�����������u8Ph4�h��,P�(h��9�����_^�M�3�賾����]ÍI W�����h�  Q�P���j�����h�R���o�������t��u��33����$    ������������@��u퍅����PhЁ������W�������������O�GG��u�f�́������f�H�H@��u���������ā�H�P������H��$    �H@��u��������j�Pj ������P�L����u/�5,Ph4�h���֋=(P��j h4�������Q��P��_^�M�3��~�����]�����������������������������������������������������������������������������������������������������������������������������������������������U���������h`�P�T��t]��3�]�������������U����   SVW��@����0   ������E�8 t��E�Q�p��B��у�;��|����E�     _^[���   ;��c�����]�������������������������������U����   SVW��@����0   �������hﾭޡp��H��@  �҃�;�����_^[���   ;��������]������������������������������U����   SVW��@����0   ������} t!��EP�p��Q��@  �Ѓ�;�����_^[���   ;��|�����]������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�p��B��  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   ������p��H��   ��;��J���_^[���   ;��:�����]����������������������U����   SVW��@����0   ������} t�E�x��u�   �3�_^[��]��������������������U����   SVW��<����1   ������=p� ��   �E��tK�}sǅ<���   �	�E��<�����MQ�UR��<���P�p��Q���   �Ѓ�;��W����\�I�}sǅ<���   �	�E��<�����MQ�UR��<���P�p��Q���  �Ѓ�;�������EP�MQ�[   ��_^[���   ;��������]���������������������������������������������������������������������U����   SVW��4����3   ������}s�E   �E��P��������E��}� u3��<�E��t�E��Pj �M�Q�������E�� �����E����E���   �E�_^[���   ;�������]������������������������������������������U����   SVW��4����3   ������} tF�E�E��=� t�E�x��u�E��P���������E�P�p��Q��Ѓ�;��w���_^[���   ;��g�����]�����������������������������������U����   SVW��@����0   ������E�p��p�� _^[��]�����������������������������U���  SVWQ�������B   ������Y�M��E��8 u3��~�E��HQ�U��BP�M��QR�E��HQ�U��
������E�}� u3��K�����$����������Pjd�����P�M��	�����Pjd�M��`���������P����������E����E�_^[��  ;��4�����]����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��E�X�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   ��Ѓ�;��N���_^[���   ;��>�����]��������������������������U���  SVWQ�������B   ������Y�M��E��8 u3���   �M�������E�M�访���E������Eԃ}� tj j�E�P�M�Q�M�载����t�E�P�ӷ����3��   �E��������tj j�M�賳���E���P�M��Qj j �U��B�M��Q�D�P�M��Q�E��H�T
�R�E��HQ�U��BP�M�Q�U��
�t��������$�������S���������Pjd�M����������������E�R��P�D蝺��XZ_^[��  ;��������]Ð   L����   Xres ����������������������������������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��E��8 u�E��@�u�����$�������L���������Pjd�����Q�U��
�������y����]荍��������������������E��H�M��E���������D{�E��u������E܋E�_^[��  ;�������]�����������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   �B<�Ѓ�;��-���_^[���   ;�������]�������������������������U���  SVWQ�������F   ������Y�M��E��8 u�E��@�u�����$�����������������Pjd�����Q�U��
�4����������]荍������������������E��H�M��E���������D{�E��u�購���E܋E�_^[��  ;��I�����]�����������������������������������������������������U����   SVW��@����0   ������p��H���   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������E�Q�p��B���   �у�;��p����E�     _^[���   ;��W�����]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q���   �Ѓ�;������_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B���   �у�;��y���_^[���   ;��i�����]� ����������������������������������U����   SVW��@����0   ������p��H����;�����_^[���   ;��������]��������������������������U����   SVW��@����0   �������E�Q�p��B�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q�p��B�H�у�;��#����E�     _^[���   ;��
�����]��������������������������������������U����   SVWQ������<   ������Y�M���h�  �E�P�� ���Q�p��B���   �у�;�������謮��������� ����w��������_^[���   ;��c�����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   �B8�Ѓ�;������_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;�����_^[���   ;��p�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�H\�у�;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�p��H���   �҃�;��z���_^[���   ;��j�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�p��B�HX�у�;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B �Ѓ�;�耾��_^[���   ;��p�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�p��B���   �у�;������_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q�B�Ѓ�;��t���_^[���   ;��d�����]� �����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�p��B��   �у�;�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q�M��B$��;��t���_^[���   ;��d�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M���x  ��;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M���|  ��;�肻��_^[���   ;��r�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;�����_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;�蝺��_^[���   ;�荺����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;��-���_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;�轹��_^[���   ;�譹����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;��M���_^[���   ;��=�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;��ݸ��_^[���   ;��͸����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;��m���_^[���   ;��]�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����  ��;������_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�p��B�H(�у�;�耷��_^[���   ;��p�����]� �������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�p��Q�B`�Ѓ�(;�����_^[���   ;��ܶ����]�$ �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�p��B�H,�у�;��`���_^[���   ;��P�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M�������P�M�������Pj j �E�P�p��Q�B4�Ѓ� ;��ȵ��_^[���   ;�踵����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;��P���_^[���   ;��@�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;�����_^[���   ;��д����]����������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q�p��B�H4�у� ;��T���_^[���   ;��D�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H�Q@�҃�;��ٳ��_^[���   ;��ɳ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�HD�у�;��\���_^[���   ;��L�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�BL�Ѓ�;�����_^[���   ;��в����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�BL�Ѓ�;��p���_^[���   ;��`�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�BP�Ѓ�;�� ���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�HT�у�;�茱��_^[���   ;��|�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�HT�у�;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H���   �҃�;�膰��_^[���   ;��v�����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�U�R�� ���P�p��Q���   �Ѓ�;������P�M������ ��������E_^[���   ;��ׯ����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q�p����   �H�у�;��T����E�_^[���   ;��A�����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�Bh�Ѓ�;��Ю��_^[���   ;��������]����������������������������U����   SVW������9   ������j �L���Ph����0�������Ph�   ������Ph�   �h�������$�����$��� t��$����t���������
ǅ���    �����_^[���   ;��
�����]������������������������������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E��M�H�E�_^[��]� �����������������������U����   SVW��@����0   ������M�C���P�M�X���P�EP�*�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E��@%��� _^[��]����������������������������U����   SVW��4����3   ������E�E��E��8 t!j �E�������E�P�3������E��     3�u�_^[���   ;��Ы����]����������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�P������E�_^[���   ;��_�����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��������M��b����E�_^[���   ;��������]��������������������U����   SVWQ��(����6   ������Y�M��M��=����E�    �	�E���E�}�}�E�M��D�    ��E�_^[���   ;��{�����]���������������������������������������U����   SVWQ��4����3   ������Y�M��M��Ǥ���M���辢��_^[���   ;�������]�����������������������U����   SVWQ��4����3   ������Y�M��M�臝��_^[���   ;�趩����]������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@`    �E��@d    �E��@h    �E����Xp�E��@x�����E��@|   _^[��]������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t j j j�E���P�M��	�����E��     �E��x` t�E���`P�ۗ����_^[���   ;�螨����]������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 tfh���P���Ph�h�h�腜����P�d�����Ph   @j膖����P諕�����(���t�h���t�3�u�3�u��E��x` tfh���P���Ph�h�h�������P�������Ph   @j������P�<������(���t�h���t�3�u�3�u��M��
����M�踪���E�P�M���dQ�U��BxP�MQ�U���`R蚒�����M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�������E��@|��   �E��xd ��   �E���pP�M���hQ�UR舥������ux�E��@h    �E����Xph���P���Ph�h�h�������P�Ȕ����Ph   @j������P�������(���t�h���t�3�u�3�u��EP�M����e���j j j�E���P�M��	�i����U��B|�E��x|t�M�訠���E��@|��E��@x�����E��@|_^[���   ;��ߥ����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVW��<����1   ������EP�+�����;Ev�M��<����	�U��<�����<���_^[���   ;�蘤����]������������������������������������U����   SVWQ��4����3   ������Y�M��M������M�蕧��_^[���   ;��.�����]��������������������������U����   SVWQ��4����3   ������Y�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	������U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[���   ;��P�����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��} t�E�M��Ap��E��xd t�E��@h��E��x|u�   �3�_^[��]� ��������������������������������U����   SVW��@����0   ������p��H����;��^���_^[���   ;��N�����]��������������������������U����   SVW��@����0   �������E�Q�p��B�H�у�;������E�     _^[���   ;��ڡ����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q�p��B�H�у� ;��T���_^[���   ;��D�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�H�у�;��ܠ��_^[���   ;��̠����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;��`���_^[���   ;��P�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H�Q�҃�;�����_^[���   ;��ٟ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M���������M������H �G@��;��_���_^[���   ;��O�����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��e������M��[����H �GD��;��Ϟ��_^[���   ;�连����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M������xH u3��#�M��ъ�����M��Ǌ�����H �FH��;��9���_^[���   ;��)�����]�������������������������������������U����   SVWQ��4����3   ������Y�M��M��S����xL u3��/��EP�MQ�UR�M��3������M��)����H �GL��;�蝝��_^[���   ;�荝����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��M�賉���xP u����3��EP�MQ�UR�EP�M�莉�����M�脉���H �WP��;������_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M������xT u����+��EP�MQ�M���������M������H �WT��;��`���_^[���   ;��P�����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��M��s����xX u����'��EP�M��Z������M��P����H �WX��;��ě��_^[���   ;�贛����]� �����������������������������U���  SVWQ�������C   ������Y�M��} t<�M��ɇ����E�P�M��χ�����M��Ň���H �WL��;��9����M��M�迊���} t?�������D���P�M腌���������s����M��|����@@�EЃ}� t�E�P�M�Z���R��P�d;聍��XZ_^[��  ;��ƚ����]� �I    l;����   x;bc ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�p��B�H�у�;������E�_^[���   ;��	�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;�蠙���E�_^[���   ;�荙����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;��0���_^[���   ;�� �����]����������������������������U����   SVWQ��4����3   ������Y�M��M��S����x` u� }  �'��EP�M��8������M��.����H �W`��;�袘��_^[���   ;�蒘����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�譄�����M�裄���H �WH��;�����_^[���   ;�������]� ��������������������������������U����   SVWQ��(����6   ������Y�M�j�EP�`����������P�M�谈���E�M�O���;E��M�w���;E�~������3��EP�MQ�UR�EP�M���������M��փ���H �WD��;��J���_^[���   ;��:�����]� ���������������������������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��M������xP u������;��EP�MQ�UR�EP�MQ�UR�M��������M��ڂ���H �GP��;��N���_^[���   ;��>�����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��c����xT u������+��EP�MQ�M��D������M��:����H �WT��;�讕��_^[���   ;�螕����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��M��Á���xX u�'��EP�M�譁�����M�裁���H �WX��;�����_^[���   ;�������]� ��������������������������������U����   SVW�� ����8   ������M�蹑���E�P�MQ���������t�}� u�M藑���E�)�E�M��U�P�M�H�U��P�M�H�U��P�ER��P��A����XZ_^[���   ;��J�����]Ð   �A����   �Adat ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E�_^[��]�����������������������������������������U����   SVW�� ����8   ������M��9����E�P�MQ�{�������t�}� u3���M�躓��R��P�4C诅��XZ_^[���   ;��������]ÍI    <C����   HCdat ������������������������������������U����   SVWQ������<   ������Y�M��M�v����M��	�����umh���T���Ph�h�h�蹆����P蘀����Ph   @j躀����P�������(���t�h���t�3�u�3�u�3��   �E�    ��E�P�M�Q�UR�E�P�p��Q���   �Ѓ�;��ّ����u3��M�E�    �	�Eԃ��EԋE�;E�}"�EԋM��<� u��EԋM���R�M�.����͍E�P�Ɂ�����   R��P��D����XZ_^[���   ;��c�����]�    �D����   �D����   �Darr count ��������������������������������������������������������������������������������������������������U����   SVWQ������?   ������Y�M��M�|���M��)�����umh���X���Ph�h�h��ل����P�~����Ph   @j��~����P��}�����(���t�h���t�3�u�3�u�3��   �E�    ��E�P�M�Q�UR�E�P�p��Q���   �Ѓ�;��������u3��u�}� u3��k�E�    �	�Eԃ��EԋE�;E�}@�EԋM��<� t�EԋM����>�����u�ϋEԋM�������������P�M�{��믍E�P�������   R��P��F����XZ_^[���   ;��[�����]�    �F����   �F����   �Farr count ����������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������p��H��   ��;�芎��_^[���   ;��z�����]����������������������U����   SVW��@����0   �������E�Q�p��B��$  �у�;�� ����E�     _^[���   ;�������]�����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�p��B��(  �у�;�虍���E�_^[���   ;�膍����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�p��B��,  �у�;�����_^[���   ;��	�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�p��B��,  �у�;�虌�������_^[���   ;�肌����]� ���������������������������U����   SVW��@����0   ������p��H��0  ��;��*���_^[���   ;�������]����������������������U����   SVW��@����0   ������p��H��4  ��;��ʋ��_^[���   ;�躋����]����������������������U����   SVW��@����0   ������p��H��p  ��;��j���_^[���   ;��Z�����]����������������������U����   SVW��@����0   ������p��H��t  ��;��
���_^[���   ;��������]����������������������U����   SVWQ��0����4   ������Y�M��} t�M�m�����0����
ǅ0���    ��0���P�M�Q�p��B��8  �у�;��v���_^[���   ;��f�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B��<  �у�;�詉��_^[���   ;�虉����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q��@  �Ѓ�;��!���_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H��D  �҃�;�覈��_^[���   ;�薈����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B��H  �у�;��)���_^[���   ;�������]� ����������������������������������U����   SVWQ������9   ������Y�M���EP�M�Q�� ���R�p��H��L  �҃�;�裇��P�M�k����� �����u���E_^[���   ;��|�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;�������E�P�MQ�p��B�H�у�;������E�_^[���   ;��ۆ����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q��T  �Ѓ�;��m���_^[���   ;��]�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B��l  �у�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q��P  �Ѓ�;��}���_^[���   ;��m�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B��X  �у�;��	���_^[���   ;��������]� ����������������������������������U����   SVW��@����0   ������p��H��\  ��;�蚄��_^[���   ;�芄����]����������������������U����   SVW��@����0   �������E�Q�p��B��`  �у�;��0����E�     _^[���   ;�������]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�p��H��d  �҃�;�蚃��_^[���   ;�芃����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�p��H��h  �҃�;��
���_^[���   ;��������]� �����������������������������������U���  SVWQ��D����o   ������Y�M��Ts���M���E��8 u�  �EP��T����s��j h�����������P��x����s��j j���T���Q��x���R������P��s����P������Q�A}����P������R�1}����P�E���)w��������؈�K�����������u���������u���������u����x����u���������Dp����T����u����K�����t�E�P��p�����2���E�$�� ����т���� ���Pjd�M��	�y���� ���耈���E�_^[�ļ  ;��o�����]� ��������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q�B�Ѓ�;��������EPj��MQ�U�R�p��H�Q�҃�;�虀���E�_^[���   ;�膀����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�Xz�����M���E�_^[���   ;��
�����]� �������������������U����   SVWQ��4����3   ������Y�M��E�P��n����_^[���   ;������]������������������������������U����   SVWQ��(����6   ������Y�M��E��8 t�E��H���M��	�E���E�}� |��E��@    _^[��]��������������������������������������U����   SVWQ������9   ������Y�M�j�M���l���E�EP�M�Q�.k�����E�3�t�E��H���U��J�E�_^[���   ;��~����]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E��8 t�E��H���M��	�E���E�}� |��E��@    _^[��]��������������������������������������U����   SVWQ��$����7   ������Y�M�j�M��yj��Pj��i������,�����,��� t$�EP��������,�������,�����$����
ǅ$���    ��$���_^[���   ;��v}����]� �����������������������������������������������U����   SVWQ������?   ������Y�M��E��HM�M�E��H�U�����M��E��M�;H��   j�EP�M��QR�Y������EȍE�P�M���Q�U��P�M��y��P�Mh�����E��}� tW�Eׅ�u-�E��8 t%�E��HQ�U�R�E��Q��k�����E�P�l�����E��M���E��MȉH�E��H�U����E��	�E��H�M�E��M�H�E�R��P�Z��n��XZ_^[���   ;��"|����]� �I    Z����   ZisRealloc ������������������������������������������������������������������������������������������U����   SVW��(����6   ������EEk��+����E��E���}�U�}� u�}� u�E+E�E��E��E�_^[��]��������������������������������������U����   SVWQ������?   ������Y�M��E��HM�M�E��H�U�����M��E��M�;H��   j�EP�M��QR�9������EȍE�P�M���Q�U��P�M��e��P��g�����E��}� tW�Eׅ�u-�E��8 t%�E��HQ�U�R�E��Q��w�����E�P�+p�����E��M���E��MȉH�E��H�U����E��	�E��H�M�E��M�H�E�R��P�(\�l��XZ_^[���   ;��z����]� �I    0\����   <\isRealloc ������������������������������������������������������������������������������������������U����   SVW��0����4   ������EPj�qe������8�����8��� t��8����U����8�����0����
ǅ0���    ��0���_^[���   ;��y����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVW��@����0   ������E��P�MQ�UR�Sr����_^[���   ;��x����]������������������������U����   SVW��,����5   ������E� j h  h����0����su��P�EP�MQ��b����_^[���   ;��w����]���������������������������������U����   SVW��@����0   ������M�b��P�M�g��P�EP�MQ�{r����_^[���   ;��1w����]�����������������������������U����   SVW��@����0   ������E��P�MQ�UR�q����_^[���   ;���v����]������������������������U����   SVW��,����5   ������E� j h  h����0����#t��P�EP�MQ�a����_^[���   ;��Uv����]���������������������������������U����   SVW��4����3   ������E��M��E�P�r�����E�     R��P�P`�h��XZ_^[���   ;���u����]�   X`����   d`tmp ����������������������������������������U����   SVW��4����3   ������E��M��E�P��q�����E�     R��P��`��g��XZ_^[���   ;��5u����]�   �`����   atmp ����������������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��4����3   ������E��M��E�P�q�����E�     R��P��a�g��XZ_^[���   ;��Ut����]�   �a����   �atmp ����������������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;���s��_^[���   ;��s����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���   �҃�;��[s��_^[���   ;��Ks����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q��  �Ѓ�;���r��_^[���   ;���r����]����������������������������������U����   SVW��@����0   ������EP�Jl����_^[���   ;��wr����]�������������������U����   SVWQ��4����3   ������Y�M��M��_v����E�P�p��Q$�BD�Ѓ�;��r���E�_^[���   ;��r����]���������������������������������U����   SVWQ��4����3   ������Y�M��M���u����E�P�p��Q$�BD�Ѓ�;��q����EP�M�Q�p��B$�Hd�у�;��vq���E�_^[���   ;��cq����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��/u����E�P�p��Q$�BD�Ѓ�;���p����EP�M�Q�p��B$�H�у�;���p���E�_^[���   ;��p����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��t����E�P�p��Q$�BD�Ѓ�;��8p����E�P�MQ�p��B$�HL�у�;��p���E�_^[���   ;��p����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q$�BH�Ѓ�;��o���M���]��_^[���   ;��xo����]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�HL�у�;��o��_^[���   ;���n����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q$�M��B��;��n��_^[���   ;��tn����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q$�M��Bl��;��n��_^[���   ;�� n����]� �������������������������U����   SVWQ��4����3   ������Y�M��p��P$��M��Bp��;��m��_^[���   ;��m����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q$�B�Ѓ�;��0m��_^[���   ;�� m����]����������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q�p��B$�H�у�;��l��P�M�s���� ����[���E_^[���   ;��l����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H�у�;��l��_^[���   ;��l����]� �������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q�p��B$�H �у�;��k��P�M�r��������F_���E_^[���   ;��rk����]� �������������������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q�p��B$�H$�у�;���j��P�M�r��������^���E_^[���   ;���j����]� �������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M��c�����X��������^���E_^[���   ;��Fj����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q$�B(�Ѓ�;���i��_^[���   ;���i����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q$�Bh�Ѓ�;��pi��_^[���   ;��`i����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H,�у�;���h��_^[���   ;���h����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H0�у�;��|h��_^[���   ;��lh����]� �������������������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q�p��B$�Ht�у�;���g��P�M��n���� ����QV���E_^[���   ;���g����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��p��P$��M��Bx��;��eg��_^[���   ;��Ug����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H4�у�;���f��_^[���   ;���f����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H8�у�;��lf��_^[���   ;��\f����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�p��B$�HL�у�;���e���E�_^[���   ;���e����]� ����������������������������������U����   SVW������9   ������EP�M��l����EP�M�Q�p��B$�H@�у�;��ee���E�P�M�ul���M��Y���ER��P��p��W��XZ_^[���   ;��-e����]�    q����   qfn �������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H@�у�;��d���E�_^[���   ;��d����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H<�у�;��d��_^[���   ;��d����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�H<�у�;��c�������_^[���   ;��c����]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H$�QP�҃�;��c��_^[���   ;��	c����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B$�HT�у�;��b��_^[���   ;��b����]� �������������������������������������U����   SVW��@����0   ������p��H$��QX��;��-b��_^[���   ;��b����]�������������������������U����   SVW��@����0   �������EP�p��Q$�B\�Ѓ�;���a��_^[���   ;��a����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q$�B`�Ѓ�;��Da��_^[���   ;��4a����]� �����������������������������U����   SVW��@����0   ������p��H(����;���`��_^[���   ;���`����]��������������������������U����   SVW��@����0   �������E�Q�p��B(�H�у�;��s`���E�     _^[���   ;��Z`����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�p��P(�M��B��;���_��_^[���   ;���_����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��p��P(��M��B��;��e_��_^[���   ;��U_����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��B��;���^��_^[���   ;���^����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�p��P(�M��B��;��y^��_^[���   ;��i^����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B(�M��P ��;���]��_^[���   ;���]����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ�p��B(�M��P��;��z]��_^[���   ;��j]����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�p��P(�M��B$��;���\��_^[���   ;���\����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��p��P(��M��B(��;��\��_^[���   ;��u\����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P(��M��B,��;��\��_^[���   ;��\����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P(��M����   ��;��[��_^[���   ;��[����]������������������������������U����   SVWQ��4����3   ������Y�M��p��P(��M��B0��;��5[��_^[���   ;��%[����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��B4��;���Z��_^[���   ;��Z����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��BX��;��PZ��_^[���   ;��@Z����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��B\��;���Y��_^[���   ;���Y����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��B`��;��pY��_^[���   ;��`Y����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��Bd��;�� Y��_^[���   ;���X����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��Bh��;��X��_^[���   ;��X����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��Bl��;�� X��_^[���   ;��X����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��Bx��;��W��_^[���   ;��W����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M����   ��;��=W��_^[���   ;��-W����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��Bt��;���V��_^[���   ;���V����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��Bp��;��`V��_^[���   ;��PV����]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��Q����t2�M��Q�M��Q����t�U��R�M���P����tǅ0���   �
ǅ0���    ��0���_^[���   ;��U����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��H����t8�MQ�A�$�M��H����t"�UQ�B�$�M���G����tǅ0���   �
ǅ0���    ��0���_^[���   ;���T����]� ������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��cB����t2�M��Q�M��PB����t�U��R�M��=B����tǅ0���   �
ǅ0���    ��0���_^[���   ;��<T����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M��\F����t<�M���A�$�M��DF����t$�U���B�$�M��,F����tǅ0���   �
ǅ0���    ��0���_^[���   ;��{S����]� ����������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��N����tE�M��Q�M��N����t2�U��R�M��N����t�E��$P�M��~N����tǅ0���   �
ǅ0���    ��0���_^[���   ;��R����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��=����tE�M��Q�M��=����t2�U��R�M��=����t�E��$P�M��}=����tǅ0���   �
ǅ0���    ��0���_^[���   ;���Q����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��K����tE�M��Q�M���J����t2�U��0R�M���J����t�E��HP�M���J����tǅ0���   �
ǅ0���    ��0���_^[���   ;��	Q����]� ��������������������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��T����tE�M��Q�M��T����t2�U��0R�M��xT����t�E��HP�M��eT����tǅ0���   �
ǅ0���    ��0���_^[���   ;��9P����]� ��������������������������������������������������U���  SVWQ�������D   ������Y�M��E�    �E�    �E�P�M���E����u3��   �}� u)��������S��P�M�A��������� >���   �   j �\���Ph��������M��P�E�RP��V�����E��}� uj��M��P��3��Lj �E�P�M�Q�M���=����u�E�P�>����3��&j �E��P�M�Q�M�>���E�P�f>�����   R��P�L��A��XZ_^[��  ;���N����]� �   T�����   n�����   l�c len ����������������������������������������������������������������������������������������������U����   SVW��8����2   ������E���8�����<����E;�8���u�M;�<���t_h�jhh��h�h���SB����P�2<����Ph   @j�T<����P�y;�����(���t�h���t�3�u�3���M��8��P�M��=��P�EP��R����_^[���   ;��M����]������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q�B�Ѓ�;���L��_^[���   ;���L����]� �����������������������������U����   SVWQ������?   ������Y�M��M��P���E�P�M��F����uǅ���    �M���:��������$�E�P�M�E:��ǅ���   �M��:�������R��P� ���>��XZ_^[���   ;��'L����]�    �����   �str ��������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�P�M�� A����u3���E�����؋M��   R��P�Ċ� >��XZ_^[���   ;��eK����]� ��   ̊����   ؊c ��������������������������������������U����   SVWQ��4����3   ������Y�M��} ����Q�M���R��_^[���   ;���J����]� ��������������������U���  SVWQ�������B   ������Y�M�j �M�B�����E�j �`���Ph���� ���� H��P�E��RP��Q�����Eԃ}� uj��M��K��3��dj �E�P�M�Q�M�>=���E�P�M��.P����t �M�Q�U�R�M���O����tǅ����   �
ǅ����    �������E�E�P�P9�����E�R��P�`��<��XZ_^[��  ;���I����]� �   h�����   t�mem ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bd��;�� I��_^[���   ;��I����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�p��P�M��Bh��;��H��_^[���   ;��H����]� ����������������������������������U����   SVWQ������<   ������Y�M��� ���P�M�j6��P�M��(Q��������� ����6�������_^[���   ;��H����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q(�M��B8��;��G��_^[���   ;��G����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q(�M��B<��;��/G��_^[���   ;��G����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q(�M��B@��;��F��_^[���   ;��F����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q(�M��BD��;��OF��_^[���   ;��?F����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��BH��;���E��_^[���   ;���E����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B(�M��P|��;��lE��_^[���   ;��\E����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q(�M��BL��;���D��_^[���   ;���D����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B(�M����   ��;��yD��_^[���   ;��iD����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�p��P(�M��BT��;���C��_^[���   ;���C����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�p��P(�M��BP��;��~C��_^[���   ;��nC����]� �����������������������U����   SVW��@����0   ������p��H(��Q��;��C��_^[���   ;��C����]�������������������������U����   SVW��@����0   �������E�Q�p��B(�H�у�;��B���E�     _^[���   ;��B����]��������������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�p��Q(�M����   ��;��	B��_^[���   ;���A����]�( ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�p��B(�H�у�;��A��_^[���   ;��uA����]���������������������������������U����   SVW��@����0   ������p��H,��Q,��;��A��_^[���   ;��A����]�������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B4��;��@��_^[���   ;��@����]���������������������������������U����   SVW��@����0   �������E�Q�p��B,�H0�у�;��C@���E�     _^[���   ;��*@����]��������������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B8��;���?��_^[���   ;��?����]���������������������������������U����   SVWQ������<   ������Y�M������P�p��Q,�M��B<��;��M?��P�M�`F���������2���E_^[���   ;��&?����]� �������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q�p��B,�M��P@��;��>��P�M�E���� ����-���E_^[���   ;��>����]� �������������������������������������������U����   SVW��@����0   �������j j �p��H,��҃�;��'>��_^[���   ;��>����]�����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H,�Q�҃�;��=��_^[���   ;��=����]� ����������������������������������U����   SVW��@����0   �������E�Q�p��B,�H�у�;��3=���E�     _^[���   ;��=����]��������������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B��;��<��_^[���   ;��<����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B��;��E<��_^[���   ;��5<����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B��;���;��_^[���   ;���;����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B ��;��e;��_^[���   ;��U;����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B$��;���:��_^[���   ;���:����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P,��M��B(��;��:��_^[���   ;��u:����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B,�M��P��;��:��_^[���   ;���9����]� �������������������������������������U����   SVWQ������<   ������Y�M������P�p��Q,�M��B��;��9��P�M�@��������:-���E_^[���   ;��f9����]� �������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H��D  �҃�;���8��_^[���   ;���8����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H��H  �҃�;��8��_^[���   ;��{8����]�����������������������U����   SVW��@����0   �������EP�p��Q��L  �Ѓ�;��"8��_^[���   ;��8����]������������������������������U����   SVW��@����0   �������EP�MQ�p��B�H�у�;��7��_^[���   ;��7����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H�Q�҃�;��>7��_^[���   ;��.7����]��������������������������U����   SVW��@����0   �������EP�MQ�p��B�H�у�;���6��_^[���   ;���6����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H�Q�҃�;��^6��_^[���   ;��N6����]��������������������������U����   SVW��@����0   �������EP�MQ�p��B�H�у�;���5��_^[���   ;���5����]�����������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;��~5��_^[���   ;��n5����]��������������������������U����   SVW��@����0   �������EP�p��Q�B�Ѓ�;��5��_^[���   ;��5����]���������������������������������U���  SVW�������E   ������E�P�M�'���M�������uǅ����    �M��Z(���������   j�E�P��+������u*�E�P�j8������uǅ����    �M��(���������Tj�EP�+������u*�EP�f7������uǅ���    �M���'��������ǅ���   �M���'�������R��P�H��&��XZ_^[��  ;���3����]�   P�����   \�parent �����������������������������������������������������������������������������U����   SVW��@����0   �������EP�p��Q�B �Ѓ�;��53��_^[���   ;��%3����]���������������������������������U����   SVW��@����0   �������EP�MQ�p��B�H(�у�;���2��_^[���   ;��2����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�p��B��  �у�;��B2��_^[���   ;��22����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q��   �Ѓ�;���1��_^[���   ;��1����]����������������������������������U����   SVW��@����0   �������EP�p��Q��  �Ѓ�;��R1��_^[���   ;��B1����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H��  �҃�;���0��_^[���   ;���0����]�����������������������U����   SVW������9   ������� ���P�p��Q�B$�Ѓ�;��r0��P�M�7���� ����$���E_^[���   ;��K0����]���������������������������������������U����   SVW������9   ������� ���P�p��Q���  �Ѓ�;���/��P�M��6���� ����#���E_^[���   ;��/����]������������������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;��N/��_^[���   ;��>/����]��������������������������U���$  SVW�������I   ������ǅ8���    �= � t!������P� ���!����8����������������K4����8���������������������������R�M�5����8�����t��8����������@"����8�����t��8�����������#"���E_^[��$  ;��O.����]�����������������������������������������������������������U����   SVW������9   �������EP�� ���Q�p��B���  �у�;���-��P�M��4���� ����x!���E_^[���   ;��-����]��������������������������������U����   SVW��@����0   ������j�EP�/�����E_^[���   ;��B-����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;���,��_^[���   ;���,����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��k,��_^[���   ;��[,����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;���+��_^[���   ;���+����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��+��_^[���   ;��{+����]�����������������������U����   SVW��@����0   ������p��H���   ��;��*+��_^[���   ;��+����]����������������������U����   SVW��@����0   �������EP�p��Q���   �Ѓ�;���*���E�     _^[���   ;��*����]�������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q�M����;��5*��_^[���   ;��%*����]� ������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M��B��;���)��_^[���   ;��)����]���������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M����   ��;��R)��_^[���   ;��B)����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B`��;���(��_^[���   ;���(����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bd��;��p(��_^[���   ;��`(����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bh��;�� (��_^[���   ;���'����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bl��;��'��_^[���   ;��'����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bp��;�� '��_^[���   ;��'����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bt��;��&��_^[���   ;��&����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��=&��_^[���   ;��-&����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M���  ��;���%��_^[���   ;��%����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bx��;��`%��_^[���   ;��P%����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;���$��_^[���   ;���$����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B|��;��$��_^[���   ;��p$����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��$��_^[���   ;���#����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��#��_^[���   ;��#����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��-#��_^[���   ;��#����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��"��_^[���   ;��"����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��M"��_^[���   ;��="����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;���!��_^[���   ;���!����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��m!��_^[���   ;��]!����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��� ��_^[���   ;��� ����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;�� ��_^[���   ;��} ����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;�� ��_^[���   ;�� ����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B��  �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M���  ��;��-��_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M����   ��;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M����   ��;��9��_^[���   ;��)����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q�p��B �H$�у�;��F����tǅ0���   �
ǅ0���    ��0���_^[���   ;������]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR�p��H �QL�҃�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q�p��B �H(�у�;�����   _^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q�M��B��;����_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q�M��B��;����_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q�M��B��;����_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M����EP�p��Q�M��B��;��?��_^[���   ;��/����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B��;��`��_^[���   ;��P����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M��P\��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M���  ��;��i��_^[���   ;��Y����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�p��P�M��B ��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$�p��P�M��B$��;��n��_^[���   ;��^����]� �����������������������U����   SVWQ��4����3   ������Y�M�����E�$�p��P�M��B(��;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B,��;����_^[���   ;��p����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B0��;����_^[���   ;�� ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B4��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B8��;��0��_^[���   ;�� ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B<��;�����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��B@��;��P��_^[���   ;��@����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��BD��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��BH��;��p��_^[���   ;��`����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��BL��;�� ��_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��BP��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q�M����   ��;����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��BT��;����_^[���   ;������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B��  �у�;��)��_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M���  ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q�M����   ��;��1��_^[���   ;��!����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q�M����   ��;����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M��PX��;��<��_^[���   ;��,����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M����   ��;�����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��M��_^[���   ;��=����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��m��_^[���   ;��]����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M����   ��;����_^[���   ;��r����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M����   ��;��	��_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M����   ��;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M���   ��;��"��_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M����   ��;��
��_^[���   ;��
����]������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M����   ��;��B
��_^[���   ;��2
����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M���  ��;���	��_^[���   ;��	����]� ����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�p��B���   �у�;��R	��_^[���   ;��B	����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q��   �Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��(����6   �������EP�MQ��,���R�p��H���  �҃�;��X��P�M� ����,��������E_^[���   ;��1����]���������������������������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;����_^[���   ;������]��������������������������U����   SVW��4����3   ������E��M��E�P�������E�     R��P��������XZ_^[���   ;��5����]�   ������   �tmp ����������������������������������������U����   SVW��@����0   ������E���Ex��M�U;�����EE�E��_^[���   ;������]� �����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B8�HD�у�;��<��_^[���   ;��,����]� �������������������������������������U����   SVW��@����0   ������p��H8��Q<��;�����_^[���   ;������]�������������������������U����   SVW��@����0   �������E�Q�p��B8�H@�у�;��c���E�     _^[���   ;��J����]��������������������������������������U����   SVW��@����0   ������p��H8����;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������E�Q�p��B8�H�у�;�����E�     _^[���   ;��j����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q8�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H8�Q�҃�;��y��_^[���   ;��i����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q8�B�Ѓ�;�� ��_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B8�H �у�;����_^[���   ;��|����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�p��H8�Q$�҃�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P�p��Q8�B�Ѓ�;��h��_^[���   ;��X����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H8�Q(�҃�;��� ��_^[���   ;��� ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q8�B,�Ѓ�;��d ��_^[���   ;��T ����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q8�B�Ѓ�;������_^[���   ;��������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R�p��H8�Q�҃�;��]���_^[���   ;��M�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H8�Q0�҃�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P�p��Q8�B4�Ѓ�;��T���_^[���   ;��D�����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B8�H8�у�;������_^[���   ;��������]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q��x  �Ѓ�;��V���_^[���   ;��F�����]����������������������������������U����   SVW��@����0   �������EP�MQ�p��B��|  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;��n���_^[���   ;��^�����]��������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�p��Q�B,�Ѓ�;��%���_^[���   ;�������]���������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP�p��Q���  �Ѓ�;�����_^[���   ;�������]��������������������������������������U����   SVW��(����6   ������M��d�����E�P�p��Q�B8�Ѓ�;������E�P�M�� ���M��u����ER��P�@�����XZ_^[���   ;��������]�   H�����   T�str ����������������������������������������U����   SVW��@����0   ������p��H��Q<��;��m���_^[���   ;��]�����]�������������������������U����   SVW��@����0   �������EP�MQ�p��B�H@�у�;�����_^[���   ;��������]�����������������������������U����   SVW��@����0   ������p��H��QD��;�����_^[���   ;�������]�������������������������U����   SVW��@����0   ������p��H��QH��;��=���_^[���   ;��-�����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H�QL�҃�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�p��B�HP�у�;��a���_^[���   ;��Q�����]�����������������������������U����   SVW��@����0   �������EP�p��Q��<  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�p��Q��,  �Ѓ�;�����_^[���   ;��r�����]������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP�p��Q���   �Ѓ�;������_^[���   ;��������]���������������������������������������U����   SVW��@����0   ������p��H�􋑼   ��;��z���_^[���   ;��j�����]����������������������U����   SVW��@����0   ������p��H���  ��;�����_^[���   ;��
�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�:  �p��B���   �у�;�����_^[���   ;�������]�����������������������������������������U����   SVW��@����0   �������EP�p��Q�B�Ѓ�;��%���_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP�p��Q��\  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW������<   ������EPj h����������P�M�Q������������������E�P�p��Q�B�Ѓ�;������M��{���R��P�8�����XZ_^[���   ;��������]Ð   @�����   L�s ��������������������������������������������������U����   SVW��(����6   ������EP�M��H����EP�M������E�P�M�0����M�������ER��P��������XZ_^[���   ;��3�����]Ë�   ������   �s ��������������������������������������U����   SVWQ��4����3   ������Y�M�j�j��EP�M��x���P�M�������E�_^[���   ;�������]� ���������������������������U����   SVWQ��4����3   ������Y�M��p��P��M��B<��;��E���_^[���   ;��5�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�p��Q�M��BL��;������_^[���   ;�������]� �����������������������������U����   SVW��@����0   �������EP�p��Q�BT�Ѓ�;��U���_^[���   ;��E�����]���������������������������������U����   SVW��@����0   �������EP�p��Q�BX�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP�p��Q�B\�Ѓ�;��u���_^[���   ;��e�����]���������������������������������U����   SVW��@����0   ������p��H��Q`��;�����_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   ������p��H��Qd��;��=���_^[���   ;��-�����]�������������������������U����   SVW��@����0   ������p��H��Qh��;������_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP�p��Q�Bl�Ѓ�;��u���_^[���   ;��e�����]���������������������������������U����   SVW��@����0   �������EP�p��Q�Bp�Ѓ�;�����_^[���   ;��������]���������������������������������U����   SVW��@����0   ������p��H���  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��2���_^[���   ;��"�����]������������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��R���_^[���   ;��B�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H�Qt�҃�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�p��Q��D  �Ѓ�;��r���_^[���   ;��b�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q��  �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������EP�MQ�p��B�Hx�у�;�����_^[���   ;��q�����]�����������������������������U����   SVW��@����0   �������EP�MQ�p��B��@  �у�;�����_^[���   ;��������]��������������������������U����   SVW������9   ������M��B�����E�P�MQ�p��B�H|�у�;������E�P�M�����M��F����ER��P�������XZ_^[���   ;��a�����]�   ������   ��fn �����������������������������������������������������U����   SVW��@����0   �������EP�MQ�p��B���   �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�p��B��h  �у�;��^���_^[���   ;��N�����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR�p��H���  �҃�;������_^[���   ;��������]���������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��k���_^[���   ;��[�����]�����������������������U����   SVW��@����0   ������p��H�􋑄   ��;��
���_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ�p��B��l  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�p��Q��   �Ѓ�;��2���_^[���   ;��"�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H��  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   ������p��H���  ��;��Z���_^[���   ;��J�����]����������������������U����   SVW��$����7   ������M��t�����E�P�p��Q���   �Ѓ�;�������E�P�M�&����M��i����ER��P�t��m���XZ_^[���   ;�������]Ð   |�����   ��bc �����������������������������������������������������U����   SVW��@����0   ������p��H��`  ��;��*���_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�p��Q��  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW�� ����8   �������EP��$���Q�p��B���   �у�;��K����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;�������]�����������������������������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP���E�$���E�$�MQ�p��B���   �у�;�����_^[���   ;�������]����������������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���   �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���   �҃�;��+���_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��K���_^[���   ;��;�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���   �҃�;��k���_^[���   ;��[�����]�����������������������U����   SVW��@����0   �������EP�MQ�p��B���   �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ�p��B���   �у�;�����_^[���   ;��~�����]��������������������������U����   SVW��@����0   �������EP�p��Q���   �Ѓ�;��"���_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�p��Q���   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�p��Q���   �Ѓ�;��B���_^[���   ;��2�����]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P�p��Q���   �Ѓ�;��������u3���E�R��P����P���XZ_^[���   ;�������]�   ������   ������   ������   ��data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P�p��Q���   �Ѓ�;��������u3���E�R��P����`���XZ_^[���   ;�������]�   ������   ������   ������   ��data sub_id main_id ������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P�p��Q���   �Ѓ�;��������u3���E�R��P�p��p���XZ_^[���   ;�������]�   x�����   ������   ������   ��data sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP�p��Q��8  �Ѓ�;�����_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�A���P�U�R�p��H0���   �҃�(;��e���_^[���   ;��U�����]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�%���P�U�R�p��H0���   �҃�(;�����_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�p��Q0���   �Ѓ�(;������_^[���   ;�������]�$ ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�p��B0���   �у�;��=���_^[���   ;��-�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q0���   �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R�p��H0���   �҃�;��F���_^[���   ;��6�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q�p��B0���   �у�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p��Q0���   �Ѓ�;��=���_^[���   ;��-�����]�������������������������U����   SVW��@����0   ������p��H0�􋑤   ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������E�Q�p��B0���   �у�;��p����E�     _^[���   ;��W�����]�����������������������������������U����   SVW��@����0   �������EP�p��Q��H  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�p��Q��T  �Ѓ�;�����_^[���   ;��r�����]������������������������������U����   SVW��@����0   ������p��H��p  ��;�����_^[���   ;��
�����]����������������������U����   SVW��@����0   ������p��H���  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��R���_^[���   ;��B�����]������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��r���_^[���   ;��b�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q���  �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW������9   �������EP�MQ�� ���R�p��H���  �҃�;��x���P�M������ ����%����E_^[���   ;��Q�����]���������������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�p��B���  �у�;������_^[���   ;��������]������������������������������U����   SVW��(����6   �������EP�MQ�UR��,���P�p��Q��X  �Ѓ�;��S���P�M�m�����,����=����E_^[���   ;��,�����]����������������������������������������U����   SVW��(����6   �������EP��,���Q�p��B���  �у�;�����P�M������,��������E_^[���   ;�������]��������������������������������U����   SVW������=   ������j hLGOg����������PhicMC�E�P�˻���������跼���M�������u�M�y����M������E��M�����P�M�:����M�������ER��P�`	聿��XZ_^[���   ;��������]Ð   h	����   t	dat ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   �BT�Ѓ�;��-���_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP�MQ�p��B��  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�p��Q��\  �Ѓ�;��R���_^[���   ;��B�����]������������������������������U����   SVW������9   ������EP��MQ�� ���R�p��H��t  �҃�;��������������� ���臾���E_^[���   ;�������]�������������������������������U����   SVW��(����6   �������EP��,���Q�p��B���  �у�;��K���P�M������,���裸���E_^[���   ;��$�����]��������������������������������U����   SVW��(����6   �������EP��,���Q�p��B���  �у�;�����P�M������,��������E_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��2���_^[���   ;��"�����]������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��R���_^[���   ;��B�����]������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ�p��B���  �у� ;������_^[���   ;�������]����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�p��H���  �҃�$;��3���_^[���   ;��#�����]�������������������������������U����   SVW��(����6   �������j �EP�MQ�UR�EP��,���Q�p��B��t  �у�;�����P�M�u�����,��������E_^[���   ;�������]����������������������������������U����   SVW��(����6   �������EP�MQ�UR�EP��,���Q�p��B���  �у�;�����P�M�)�����,���������E_^[���   ;��������]������������������������������������U����   SVW��@����0   �������EP�p��Q��8  �Ѓ�;�����_^[���   ;��r�����]������������������������������U����  SVW��(����6  �����󫡐�3ŉE��E�E�E�P�MQh   ������R�T�����������Ph��p��Q��4  �Ѓ�;�������E�    R��P�|�q���XZ_^[�M�3�贰�����  ;�������]ÍI    �����   �t ��������������������������������������������������������������U����   SVW��4����3   ������} 3��   �EP�MQ�UR�EP�������E��}� |�E��9E�|�}� }fh��d���Ph�h�h��3�����P������Ph   @j�4�����P�Y������(���t�h���t�3�u�3�u��EE�@� �E���E��E�_^[���   ;��h�����]��������������������������������������������������������������������U����   SVW��(����6   �������,���P�p��Q��  �Ѓ�;������P�M������,����7����E_^[���   ;�������]������������������������������������U����   SVW��(����6   �������,���P�p��Q��  �Ѓ�;��O���P�M������,���觰���E_^[���   ;��(�����]������������������������������������U����   SVW������=   ������������u�\h���M��^����EPh���M��2����EPh���M��!���j �E�PhicMC�����Q�+���������������M�����R��P������XZ_^[���   ;��[�����]Ë�   �����   �msg ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�p��B�M��P4��;�����_^[���   ;�������]� �������������������������������������U����   SVW������=   ������聬����u�M�{����E�^h!���M��Ӵ���EPh!���M�觶��j �E�PhicMC�����Q豮�������V���P�M����������������M�腯���ER��P�X色��XZ_^[���   ;��ο����]Ð   `����   lmsg ����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   �BH�Ѓ�;��-���_^[���   ;�������]�������������������������U����   SVW������=   ������������u�M������E�^h����M��S����EPh����M��'���j �E�PhicMC�����Q�1��������֭��P�M�V���������x����M������ER��P���	���XZ_^[���   ;��N�����]Ð   �����   �msg ����������������������������������������������������������������U���   SVW�� ����@   ������������u3��^h#���M��L����EPh#���M�� ���j �E�PhicMC�����Q�*�������詪�������������t����M����������R��P������XZ_^[��   ;��G�����]Ë�   �����   �msg ��������������������������������������������������������U���   SVW�� ����@   ������������u3��^hs���M��L����EPhs���M�� ���j �E�PhicMC�����Q�*�������詩�������������t����M����������R��P������XZ_^[��   ;��G�����]Ë�   �����   �msg ��������������������������������������������������������U����   SVW��@����0   ������p��H��d  ��;�躻��_^[���   ;�誻����]����������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP�p��Q��h  �Ѓ�;��:���_^[���   ;��*�����]��������������������������������������U����   SVW��@����0   �������EP�MQ�p��B��l  �у�;�辺��_^[���   ;�论����]��������������������������U����   SVW��@����0   ������p��H�􋑄  ��;��Z���_^[���   ;��J�����]����������������������U����   SVW��$����7   �������EP��(���Q�p��B���  �у�;�����P�M�*�����(����j����E_^[���   ;��Ĺ����]��������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��b���_^[���   ;��R�����]������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�p��B���  �у�;��~���_^[���   ;��n�����]��������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;�蛷��_^[���   ;�苷����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��+���_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H��l  �҃�;�軶��_^[���   ;�諶����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��K���_^[���   ;��;�����]�����������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;�����_^[���   ;��ҵ����]������������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��r���_^[���   ;��b�����]������������������������������U����   SVW��@����0   �������EP�MQ�p��B��$  �у�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�p��Q��(  �Ѓ�;�蒴��_^[���   ;�肴����]������������������������������U����   SVW��@����0   �������EP�p��Q��,  �Ѓ�;��"���_^[���   ;�������]������������������������������U����   SVW��@����0   ������p��H��0  ��;�躳��_^[���   ;�誳����]����������������������U����   SVW��@����0   ������p��H��<  ��;��Z���_^[���   ;��J�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�p��Q���  �Ѓ�;�����_^[���   ;��ֲ����]����������������������������������U����   SVW��@����0   ������p��H���  ��;��z���_^[���   ;��j�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;�����_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�p��Q��   �Ѓ�;�袱��_^[���   ;�蒱����]������������������������������U����   SVW��4����3   ������j �M�����E��}� t�E�P��������E�P茠����R��P� %�£��XZ_^[���   ;�������]Ë�   (%����   4%c ������������������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ�p��B��  �у� ;��f���_^[���   ;��V�����]����������������������������������U����   SVW��@����0   ������p��H��P  ��;������_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H��`  �҃�;�苯��_^[���   ;��{�����]�����������������������U����   SVWQ��4����3   ������Y�M��E���P�g�����_^[���   ;�������]���������������������������U����   SVW��@����0   �������EP�p����   ���   �Ѓ�;�迮��_^[���   ;�诮����]���������������������������U����   SVW��@����0   ������jjj������P�ڜ����P�EP�8�Q�C�����P�:�������u�   j�EP�#�������th ��_������j�EP��������th��>������EP�2�����h   @�EP�ԗ������t�EP�MQ�'  ��h    �EP诗������uh�������_^[���   ;�蓭����]�������������������������������������������������������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVW��@����0   ������EPh�蓭����_^[���   ;��¬����]������������������������������U���0  SVW�������L  �����󫡐�3ŉE��E�P�o  ���E�P�  ���E�E�Ph<�j?�M�Q�~������EP�MQ�U�Rh,�h�  ������P謘����������P�[�����R��P�@*譞��XZ_^[�M�3�������0  ;�������]ÍI    H*����   {*����@   p*����   l*dst timestring rawtime �����������������������������������������������������������������������������U����   SVW��@����0   ������EP�0�����_^[���   ;�������]�������������������U����   SVW��@����0   ������EP臭����_^[���   ;��Ǫ����]�������������������U����   SVW��(����6   ������} 3��   �E�E��E�P�MQ�UR�EP�_������E�}� |�E�;E|�}� }fhH��l���Ph�h�h�萞����P�o�����Ph   @j葘����P趗�����(���t�h���t�3�u�3�u��EE�@� �E���E��E�    �E�_^[���   ;�辩����]��������������������������������������������������������������������������U����  SVW��(����6  �����󫡐�3ŉE�h    �8�P�1�������t
耗���8�jjj蘗����P菗����P�EP�8�Q�������P��������u��   �E������������P�MQh�  ������R�]�����j�EP谒������th ��������j�EP菒������th��ˤ����������P輤����h   @�EP�^�������t�EP�MQ������h    �EP�9�������uh��u�����ǅ����    R��P�0.轚��XZ_^[�M�3�� ������  ;��������]ÍI    8.����   D.t ����������������������������������������������������������������������������������������������������������U����   SVW��@����0   ������h    jjj辕����P赕����P謕����_^[���   ;�������]��������������������������U����   SVW��@����0   ��������X;��Ԧ�������_^[���   ;�辦����]��������������������������U����   SVWQ��4����3   ������Y�M��E�� P��E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M��g����E��t�E�P�������E�_^[���   ;��������]� ������������������������U����   SVWQ��4����3   ������Y�M��E�� P�_^[��]��������������U����   SVWQ������9   ������Y�M��E��E�E�E��E��8 t2��j �E���U����ȋ��;��M����E�P�A������E��     3�u�R��P�1�Η��XZ_^[���   ;�������]Ë�   1����   (1_this ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M���  ��;�肤��_^[���   ;��r�����]������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M���(  ��;�����_^[���   ;�������]������������������������������U����   SVWQ������<   ������Y�M������P�p��Q�M���   ��;�蚣��P�M譪��������G����E_^[���   ;��s�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��p��P��M���$  ��;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�p��B��  �у�;�莢��_^[���   ;��~�����]��������������������������U����   SVW��@����0   �������EP�p��Q���  �Ѓ�;��"���_^[���   ;�������]������������������������������U����   SVW��@����0   ������p��H��  ��;�躡��_^[���   ;�誡����]����������������������U����   SVW��@����0   �������EP�MQ�UR�p��H���  �҃�;��K���_^[���   ;��;�����]�����������������������U����   SVW��@����0   �������EP�MQ�p��B��x  �у�;��ޠ��_^[���   ;��Π����]��������������������������U����   SVW��@����0   �������EP�p��Q��|  �Ѓ�;��r���_^[���   ;��b�����]������������������������������U����   SVW��@����0   ������p��H��d  ��;��
���_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ�p��B��p  �у�;�螟��_^[���   ;�莟����]��������������������������U����   SVW��@����0   �������EP�MQ�p��B��t  �у�;��.���_^[���   ;�������]��������������������������U����   SVW��4����3   ������E��M��E�P�X������E�     R��P��7�`���XZ_^[���   ;�襞����]�   �7����   �7tmp ����������������������������������������U����   SVWQ��4����3   ������Y�M���j j��p��P�M��B��;��!����E�_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���j �EP�p��Q�M��B��;�讝���E�_^[���   ;�蛝����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���EPj��p��Q�M��B��;��.����E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M�輦��_^[���   ;�趜����]������������������U����   SVWQ��4����3   ������Y�M��p��P��M��B��;��e���_^[���   ;��U�����]���������������������������������U����   SVWQ��4����3   ������Y�M�j j �E�P�M�3����E�_^[���   ;�������]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�p��P�M����   ��;�膛��_^[���   ;��v�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�H�у�;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p��B�H�у�;�茚�������_^[���   ;��u�����]� ������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��q����E�M��ۏ��_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   �BX�Ѓ�;�蝙��_^[���   ;�荙����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M��Bt��;��0���_^[���   ;�� �����]� �������������������������U����   SVWQ��4����3   ������Y�M�h#  �EP�MQ�M�荄��_^[���   ;�蹘����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�p��P�M��Bl��;��I���_^[���   ;��9�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�hF  �EP�MQ�M�蝃��_^[���   ;��ɗ����]� ����������������������������������U����   SVWQ��(����6   ������Y�M��EP�M�������E�EP�M��˄��_^[���   ;��S�����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q�p����   �H`�у�;�����_^[���   ;��ٖ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�p��Q�M����   ��;��m���_^[���   ;��]�����]� ����������������������U����   SVWQ��(����6   ������Y�M���EP�p��Q�M����   ��;�������E�}� u3���M�����_^[���   ;��ؕ����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P�p����   �B�Ѓ�;��m���_^[���   ;��]�����]�������������������������U����   SVW��4����3   ������j�   ���E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;��Ҕ��_^[���   ;������]����������������������������������������������U����   SVW��@����0   ������h��EPh�f ������_^[���   ;��M�����]�������������������������U����   SVW������<   ������j�{������E��}� t	�E��x uǅ��������M覇��������E�E8P�M4Q�U0R�E,P�M(Q���̍UR�ך���EP�M��Q�҃�4�� ����M�_����� ���_^[���   ;�舓����]����������������������������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;������_^[���   ;�������]�����������������������������������U����   SVW��4����3   ������j�������E��}� t	�E��x u3����EP�M��Q�҃�;��k���_^[���   ;��[�����]���������������������������������������U����   SVWQ������>   ������Y�M���EP�p��Q�M��Bd��;������E�}� u3��nj �����Phd�������u���P�E���RP� ������E��}� u3��4��EP�M��Q�U�R�p��P�M��Bh��;�聑���E�E��  �E�_^[���   ;��e�����]� ��������������������������������������������������������������U����   SVW��@����0   ������j h�  h`��M�����`�_^[���   ;��ڐ����]����������������������U����   SVW��@����0   ������j h�  h`��M蒃���`�_^[���   ;��z�����]����������������������U����   SVW��@����0   ������h� �M辅����tj h�  h`��M� ����������h��h`��Є�����`�_^[���   ;�������]������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�p����   �M��B��;��}���_^[���   ;��m�����]� ����������������������U����   SVWQ��4����3   ������Y�M��p����   ��M��Bx��;�����_^[���   ;�������]������������������������������U����   SVW��(����6   ������j h�  h`���,���P�M��|����褁����,����}���`�_^[���   ;�聎����]�����������������������������U����   SVW��(����6   ������j h�  h`���,���P�M�S|�����$�����,����|���`�_^[���   ;�������]�����������������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ��w����_^[���   ;�萍����]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��(����6   ������j�EP��������E��}� u3���M������E�3��}� ��_^[���   ;��Ԍ����]��������������������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�g������E��}� u3��5�M��W����E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;�������]���������������������������������������%L�%P�%T�%X�%(�%,U��W�}3�������ك��E���8t3�����_��������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �E�����3��} ���E��}� uh�j j.hx�j�|������u̃}� u+�����    j j.hx�hd�h�����������W�U�B��@t�M�A    �=�UR�v������E�    �EP�v�����E��E������   ��MQ�i�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������̋�U����E�����3��} ���E�}� uh8�j jYhx�j�[{������u̃}� u.輒���    j jYhx�h�h8��ǌ��������   �U�U��E��H��   ta�U�R�F������E��E�P�~�����M�Q� �����P�ȏ������}	�E������$�U��z tj�E��HQ�������U��B    �E��@    �E���]�����������������������������������������������������������������������̋�U��Q�E�    �} u3��S  �}��   �	�E����E��M��9M���   �U���U�E���E�M�Q���t�E�H��U�B�;�t�M�A��U�J�+���   �U�B���t�M�Q��E�H�;�t�U�B��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��   �E�H���t�U�B��M�Q�;�t�E�@��M�Q�+��X�����	�E����E��M�;Ms>�U���t�M��E�;�t�U��M�+���E���E�M���M�3���]�����������������������������������������������������������������������������������������������̋�U��j�h�h9�d�    P�ĸSVW���1E�3�P�E�d�    �E�E܋M�M��} u�} t	�E�    ��E�   �U��Uԃ}� uh`�j j7h��j�x������u̃}� u-�g����    j j7h��h��h`��r�����3���  3Ƀ} ���MЃ}� uh��j j8h��j�w������u̃}� u-�����    j j8h��h��h��������3��`  3��} ���Ẽ}� uh��j j9h��j�@w������u̃}� u-衎���    j j9h��h��h��謈����3���  �} u3���  �U�U�E�P�7������E�    �M�MȋUȋB��@��   �M�Q�������Eă}��t!�}��t�U����Eă�������E���E����M��Q$������uA�}��t!�}��t�M����Uă�������U���E����E��H$�� ���х�t	�E�    ��E�   �E��E��}� uh`�j jJh��j�	v������u̃}� u-�j����    j jJh��h��h`��u������E�    �}� ��   �U���U��   �E�H���M��U�E��B�}� |�M��%�   �E��M����E���M�Q��}�����E��U��U؃}��u�E�;Eu	�E�    �)�!�M܊U؈�E؋M܃��M܃�
u��h����U�� �E������   ��E�P者����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    3��} ���E܃}� uh��j j6h �j�s������u̃}� u-�����    j j6h �h�h��������3��V  3҃} �U؃}� uh�j j7h �j�Gs������u̃}� u-訊���    j j7h �h�h�賄����3���   �M�����ډU�uh��j j8h �j��r������u̃}� u-�F����    j j8h �h�h���Q�����3��   誊���E�}� u�����    3��t�E�    �M���u*�����    �E�    j��E�Ph���s�����E��9�M�Q�UR�EP�MQ�z�����E��E������   ��U�R葂����ËE��M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������̋�U��j@�EP�MQ��w����]�������̋�U��Q3��} ���E��}� u!hȑj h�   h �j�1q������u̃}� u0蒈���    j h�   h �h��hȑ蚂�����   �-h�   �UR�EP�pw�����M��U�: t3���<���� ��]������������������������������������������������̋�U��j�hH�h9�d�    P���SVW���1E�3�P�E�d�    3��} ���E؃}� uht�j j6h �j�8p������u̃}� u.虇���    j j6h �h�ht�褁��������   �U�U��|���� Pj�0������E�    �e|���� P�do�����E܋E�Pj �MQ�G|���� P�f|�����E��3|���� P�U�R茄�����E������   ��|���� Pj�����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�^h������]������������̋�U��Q�E�E��M�Q�UR�EP��s������]������������̋�U��Q�E�E��M�Qj �UR�s������]��������������̋�U��Q�E�E��M�Q�UR�EP�s������]������������̋�U��Q�E�E��M�Qj �UR�qs������]��������������̋�U��������3�9�����M��} t������U���E�    �E�����E���]������������������������̋�U�졐���3�9������]��������������������̋L$W����   VS�ًt$��   �|$u����   �'��������t+��t/��   u����ua��t��������t7��u�D$[^_���   t�������   ��   u����ut�����u�[^�D$_É����t�����~�Ѓ��3��� �t܄�t,��t��  � t��   �uĉ�����  �����   ��3҉��3���t3������u����w����D$[^_�����������������������������������������������������������������������������;��u���
n������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    �}��   �f����u3��  �u����u�o��3��  �z���p�	�]�������;y����}�nt���Ko��3��i  蝄����|辂����|j �^�������t��q���8t���o��3��3  j��������������  �} um�=�� ~X���������E�    �=� u�j���lq����s���n���E������   ��} u�=��t�s����3��   �   �}��   ��c��h�   h��jh  j�������E�}� tV�U�R��P���Q�l�Ѕ�t%j �U�R��~�����h�M��U��B�����j�E�P�Ox����3���3����}u
j �9m�����   �M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��}u�h���EP�MQ�UR�   ��]� �����������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �e��E�   �} u�=�� u3��N  �E�    �}t�}uT�=�� t�EP�MQ�UR����E�}� t�EP�MQ�UR�V���E�}� u�E�    �E������E���   �EP�MQ�UR�'e���E�}u=�}� u7�EPj �MQ�	e���URj �EP��~���=�� t�MQj �UR����} t�}u@�EP�MQ�UR��~����u�E�    �}� t�=�� t�EP�MQ�UR����E��E������8�E���U��E�P�M�Q�Lo����Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������u�U��� PRSVW�Ej P�0}����_^[ZX��]�����������̋�U��QSVW3���ى}�9>~H���$    ��F�8�|�����u�T8с<����t�L8�UQR��k�����E�@���E�;|�_^[��]���������������������������̋�U��V���t!��tS�]��tW�̋�����F�V�3_[^]� �������������̋�U��QSVW��3���;�tR�}�9>~K��    �F�8�����9T�u�D8�9t�N�T�ERP�k��������̋E�@���E�;|������̋u3��ƅ�tV�@G��u���tJ9u9Vu
9Vu9Vt�MWVQ�2|��������̋F9T0�t�MWVQ�|��������̋vO��u�_^[��]� �����������������������������������������������������������̀=�� uj jj j j ����w��P�Jn����������������������������jjj j j �lw�����������������̋T$�L$��ti3��D$��u���   r�=<� t�^k��W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$��������������������������������������̋�U��Qj j j���P�MQ��r�����E��E���]������������������������̋�U��j�EP��q����]�����������̋�U���_m���} t�=\����]�������̋�U���0�C��4����8�_��<�^��@����D�C��H����L� ��P���T���]�������������������������������������̋�U��Q����E��M����E���]������������������̃=<� t-U�������$�,$�Ã=<� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������������������������������������������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+���������������������������������������U��WV�u�M�}�����;�v;���  ���   r�=<� tWV����;�^_u��]����   u������r)��$��g�Ǻ   ��r����$��f�$��g��$�Tg��fg4g#ъ��F�G�F���G������r���$��g�I #ъ��F���G������r���$��g�#ъ���������r���$��g�I �g�g�g�g�g�g|gtg�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��g���g�g�g�g�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�\i�����$�i�I �Ǻ   ��r��+��$�`h�$�\i�ph�h�h�F#шG��������r�����$�\i�I �F#шG�F���G������r�����$�\i��F#шG�F�G�F���G�������V�������$�\i�I ii i(i0i8i@iSi�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�\i��liti�i�i�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���(V�E�    �EP�M��f���M��1\������   �U��E�    �	�E����E��}�s3�M��U��P�_�������M��U�D�P�_����E��L0�M��jXhx�j�U���R�?V�����E��}� ��   �E��E��E�    �	�M����M��}���   �U��:�E܃��E�j j_h �h�hh��M��U��P�M����U�+U�+�Q�E�P�dt����P�f�����M�Q��^����E܉E܋U��:�E܃��E�j jbh �h�h���M��U�D�P�M����U�+U�+�Q�E�P�t����P�Bf�����M�Q�u^����E܉E��#����U�� �E܃��E܋M��M؍M��:s���E�^��]����������������������������������������������������������������������������������������������������������������̋�U��} u��EP�MQ�UR�EP�MQ��k��]������������������������̋�U��Q�M��E��@ �} ��   �b���M��A�U��B�M��Pl��E��H�U��Ah�B�M��;D�t�E��H�Qp#��u
�i���M���U��B;��t�M��Q�Bp#��u�#k���M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������������������������������������������������������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]�������������������̋�U��Q�M��E���]����������������̋�U��j ��n����]���������������̋�U���(V�E�    �EP�M��b���M��AX������   �U��E�    �	�E����E��}�s4�M��U�D�8P�[�������M��U�D�hP�[����E��L0�M��jhx�j�U���R�NR�����E��}� �  �E��E��E�    �	�M����M��}���   �U��:�E܃��E�j h�   h �h��h(��M��U�D�8P�M����U�+U�+�Q�E�P�op����P�b�����M�Q��Z����E܉E܋U��:�E܃��E�j h�   h �h��h���M��U�D�hP�M����U�+U�+�Q�E�P�	p����P�Jb�����M�Q�}Z����E܉E������U�� �E܃��E܋M��M؍M��Bo���E�^��]������������������������������������������������������������������������������������������������������������������������̋�U��j �a����]���������������̋�U���,V�E�    �EP�M��g`���M���U������   �U��E�    �	�E����E��}�s3�M��U��P�\Y�������M��U�D�P�GY����E��L0�M���E�    �	�U����U��}�s4�E��M�T�8R�Y�������E��M�T�hR��X����E��D0�E�뽋M􋑘   R��X�������E􋈜   Q��X����E��T0�U��E􋈠   Q�X�����U��D�E��M􋑤   R�X�����M��T�U��E􋈨   Q�uX�����U��D�E��M���d  �M�h�   hx�j�U�R�#O�����E��}� ��  �E��E؋M���d  �M�hd  �U�R�E�P�b^�����E�    �	�M����M��}���   �U��E؋M܉�j h�   h �ht�h��U��E��Q�U�+U��E�+�P�M�Q�*m����P�k_�����U�R�W�����M܍T�U܋E��M؋U܉T�j h�   h �ht�h���E��M�T�R�E�+E��M�+�Q�U�R��l����P�_�����E�P�9W�����M܍T�U�� ����E�    �	�E����E��}���   �M��U؋E܉D�8j h�   h �ht�h8��M��U�D�8P�M�+M��U�+�R�E�P�?l����P�^�����M�Q�V�����U܍D�E܋M��U؋E܉D�hj h�   h �ht�hЗ�M��U�D�hP�M�+M��U�+�R�E�P��k����P�^�����M�Q�NV�����U܍D�E������M؋U܉��   j h�   h �ht�hp��E􋈘   Q�U�+U��E�+�P�M�Q�rk����P�]�����U�R��U�����M܍T�U܋E؋M܉��   j h�   h �ht�h��U􋂜   P�M�+M��U�+�R�E�P�k����P�P]�����M�Q�U�����U܍D�E܋M؋U܉��   j h�   h �ht�h���E􋈠   Q�U�+U��E�+�P�M�Q�j����P��\�����U�R� U�����M܍T�U܋E؋M܉��   j h�   h �ht�h0��U􋂤   P�M�+M��U�+�R�E�P�Ij����P�\�����M�Q�T�����U܍D�E܋M؋U܉��   j h�   h �ht�hȕ�E􋈨   Q�U�+U��E�+�P�M�Q��i����P�'\�����U��UԍM��Ei���E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �
M����]���������������̋�U��EPj �MQ�UR�EP�MQ�nK����]�����������̋�U��j j �EP�MQ�UR�EP�@K����]�������������̋�U��j �EP�MQ�UR�EP�MQ�K����]�����������̋�U���\�E�    �E�E��MQ�M���X��3҃} �U؃}� u!h̚j hK  h �j��N������u̃}� u@�Gf���    j hK  h �h��h̚�O`�����E�    �M��f���E���  3Ƀ} ���Mԃ}� u!h��j hL  h �j�mN������u̃}� u@��e���    j hL  h �h��h����_�����E�    �M��'f���E��P  �E�  3Ƀ} ���MЃ}� u!hX�j hO  h �j��M������u̃}� u@�Oe���    j hO  h �h��hX��W_�����E�    �M��e���E���  �} u�M��M��� ���   �M���U�U��E��E܋M�M��}� ��  �U��E��}� t�}�%t
��   �  3Ƀ} ���M̃}� u!h0�j hp  h �j� M������u̃}� u@�d���    j hp  h �h��h0��^�����E�    �M���d���E��  �E���E�E�    �M���#u�E�   �E���E�M�Q�U�R�E�P�MQ�UR�E�Q�M���K��P��  ����u�}� v�E�   �   �U���U�   �M���K��P�E�Q�M������tf�}�v`�U�B��u03�u!h��j h�  h �j�L������u��E�   �Q�%�E�M���E���E�M���M�U����U��E�M���E���E�M���M�U����U��8����}� u*�}� v$�E�  �M+M��M��M��c���E��   �   �U�� �}� u�}� w��b��� "   �q�E�    �}� u!h��j h�  h �j�6K������u̃}� u=�b���    j h�  h �h��h���\�����E�    �M���b���E���E�    �M���b���E���M���b����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   V�E�E��M����M��}�v��  �U�����$����M�y |�U�z	�E�   ��E�    �E��E�}� u!h��j h  h �j�4I������u̃}� u0�`���    j h  h �hp�h���Z����3��(  �UR�EP�M�Q�E��Q��  ���  �U�z |�E�x	�E�   ��E�    �M��M��}� u!h��j h  h �j�H������u̃}� u0��_���    j h  h �hp�h����Y����3��  �EP�MQ�U�B�M�T�R�B  ���Y  �E�x |�M�y	�E�   ��E�    �U��U�}� u!h�j h   h �j��G������u̃}� u0�F_���    j h   h �hp�h��NY����3���  �MQ�UR�E�H�U�D�8P�  ���  �M�y |�U�z	�E�   ��E�    �E��E�}� u!h�j h(  h �j�=G������u̃}� u0�^���    j h(  h �hp�h��X����3��1  �UR�EP�M�Q�E�L�hQ��  ���	  �}  ��   �UR�EP�MQ�URj�EP��  ����u3���  �M�9 u3���  �U��  �M����E��M����E��MQ�UR�EP�MQj�UR�  ����u3��  �   �EP�MQ�UR�EPj �MQ�]  ����u3��S  �U�: u3��D  �E�� �U����M��U����M��UR�EP�MQ�URj�EP�  ����u3���
  ��
  �M�y|�U�z	�E�   ��E�    �E��E�}� u!hX�j hg  h �j�{E������u̃}� u0��\���    j hg  h �hp�hX���V����3��o
  �U R�EP�MQj�U�BP�  ���H
  �M�y |�U�z	�E�   ��E�    �E��E��}� u!hȝj hp  h �j��D������u̃}� u0�5\���    j hp  h �hp�hȝ�=V����3���	  �U R�EP�MQj�U�BP��  ���	  �M�y |�U�z	�E�   ��E�    �E��E܃}� u!hȝj hx  h �j�-D������u̃}� u0�[���    j hx  h �hp�hȝ�U����3��!	  �U�B��   ���U��}� u�E�   �U R�EP�MQj�U�R�(  ����  �E�x |�M�ym  	�E�   ��E�    �U��U؃}� u!h8�j h�  h �j�hC������u̃}� u0��Z���    j h�  h �hp�h8���T����3��\  �M Q�UR�EPj�M�Q��R�{  ���2  �E�x |�M�y	�E�   ��E�    �U��Uԃ}� u!h�j h�  h �j�B������u̃}� u0�Z���    j h�  h �hp�h��'T����3��  �M Q�UR�EPj�M�Q��R��  ���  �E�x |�M�y;	�E�   ��E�    �U��UЃ}� u!h��j h�  h �j�B������u̃}� u0�uY���    j h�  h �hp�h���}S����3��  �M Q�UR�EPj�M�QR�*  ����  �E�x |�M�y	�E�   ��E�    �U��Ũ}� u!hȝj h�  h �j�mA������u̃}� u0��X���    j h�  h �hp�hȝ��R����3��a  �M�y�UR�EP�M���   R�  ����EP�MQ�U���   P�  ���  �M�9 |�U�:;ǅ|���   �
ǅ|���    ��|����Eȃ}� u!h(�j h�  h �j�@������u̃}� u0��W���    j h�  h �hp�h(��R����3��  �U R�EP�MQj�U�P�
  ���k  �M�y |�U�zǅx���   �
ǅx���    ��x����Eă}� u!h��j h�  h �j��?������u̃}� u0�OW���    j h�  h �hp�h���WQ����3���  �U�B�E��a  �\  �M�y |�U�zǅt���   �
ǅt���    ��t����E��}� u!h��j h�  h �j�M?������u̃}� u0�V���    j h�  h �hp�h���P����3��A  �U R�EP�MQj�U�BP�c	  ���  �M�y |�U�zǅp���   �
ǅp���    ��p����E��}� u!h��j h�  h �j�>������u̃}� u0��U���    j h�  h �hp�h���P����3��  �U�z u	�E�   ��E�H���M��U�z |�E�xm  ǅl���   �
ǅl���    ��l����M��}� u!h8�j h�  h �j��=������u̃}� u0�OU���    j h�  h �hp�h8��WO����3���  �E�H;M�}	�E�    �-�U�B��   ���E��U�B��   ��;U�|	�U����U��E P�MQ�URj�E�P��  ���}  �}  t+�MQ�UR�EP�MQj�UR�]	  ����u3��S  �)�EP�MQ�UR�EPj �MQ�2	  ����u3��(  �  �UR�EP�MQ�URj�EP�	  ����u3���  ��  �M3҃y �U��}� u!h�j h�  h �j�<������u̃}� u0��S���    j h�  h �hp�h���M����3��  �M�A��d   ���U��U R�EP�MQj�U�R�  ���T  �E�x����|�M�y�  ǅh���   �
ǅh���    ��h����U��}� u!hX�j h  h �j��;������u̃}� u0�2S���    j h  h �hp�hX��:M����3���   �M�A��d   ���ȃ�k�d�U�B��d   ��ʉM��E P�MQ�URj�E�P��  ���{�:���MQ�UR�=���M3҃y  ��P�5  ���O�M��%�E����U�
�E����U�
�+�)3�u!h �j h  h �j��:������u�3���   ^��]ÍI t�P��~�W������4�����K�$��}F������m���Շ"���v�  	
������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�8 t;�M���t1�E��U���M����E��M���M�U����M��]����������������������̋�U��Q�E�    �} t�EP�MQ�UR�   ���}�E�M;sj�U���U�	�E���E�M��t2�E��
   ����0�E��E��E��
   ���E�U����U�뽋E�M��U�
�E�+M��U�
�	�E�     ��]������������������������������������������������������̋�U����E��M��U�:vE�E��
   ����0�E���M����M��U����M��E��
   ���E�} ~�U�:w��E��M�U�E���M����M��U���E��M��U���M����M��U�E���M���M�U�;U�r̋�]��������������������������������������������������̋�U���\���3ŉE��E�Eă}� t�}�t��M���   �U���E���   �M���U���   �E�M���   �?  �}t�x�U���t�E̋M�Q��l  f�UЋE�H��f�MҋUf�Bf�E֋Mf�Qf�U؋Ef�Hf�MڋUf�f�E�3�f�M�j j �U�R�E�Pj �M���   R�ỦE�}� ��   h��  �E��P��5����P�G�����Eȃ}� ��   �M�Q�U�R�E�P�M�Qj �U���   P�ỦE�MȉM��U���U�}� ~9�E�8 v1�M��E���
�U����M��U����U��E����U�
븋E�P�NH�����   ��  �M������  �E�8 ��  �E� �E�    �E�    �M�M��	�U����U��E���U���U����U�;�u�܋E����E��M���U��E���'�E��}�R�b  �M���T��$�(��E��E��M����M��}�w!�U��$����E�   �E�m�
�E�b��E�B�  �E��E��M����M��}�w!�U��$����E�   �E�d�
�E�a��E�A��  �E��E��}�t�}�t�
�E�y��E�Y�  �M��M��}�t�}�t	��E�   �E�I�  �U��U��}�t�}�t	��E�   �E�H�p  �E��E��}�t�}�t	��E�   �E�M�L  �M��M��}�t�}�t	��E�   �E�S�(  hT��U�R�2������u�E���E��hP��M�Q��1������u	�U���U��E�p��  �E�x�M���   �U���E���   �M��}���   �U�: ��   �EP�M��R�<1������tn�E�8vf�M��Q��u,3�u!h��j h�  h �j�/������u�3��P  �U��M����E����U�
�E����E��M����E��M��E���
�U����M��U����U��E����U�
��   �E������   �U�: ��   �EP�M��R�i0������tn�E�8vf�M��Q��u,3�u!h��j h�  h �j��.������u�3��}  �U��M����E����U�
�E����E��M����E��M��E���
�U����M��U����U��E����U�
�-����E��E��2����M�����   �U�U��U�E������   �U�: ��   �E����'u�U���U��   �EP�M��R�]/������tn�E�8vf�M��Q��u,3�u!h �j h�  h �j��-������u�3��q  �U��M���E����U�
�E���E�M����E��M��E��
�U����M��U���U�E����U�
�����	�E�E��E��!����M��t;�U�R�EP�MQ�UR�EP�M�Q�UR�z�������u3���   �E��E��   �MQ�U��P�Q.������tk�M�9vc�U��B��u)3�u!h �j h�  h �j��,������u�3��h�E��U���M����E��M���M�U����M��U��M���E����U�
�E���E�M����E��(����   �M�3���&����]������˕�d���Ж;�A�� 







































































	�������%�,�2�8��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP��?�����.�}���  t%3�u!hءj h�   h`�j�)������u̋�]��������������������������̋�U���4VW�E�    �E�    �E�    �E�    3��} ���E��}� uh��j jEh@�j�(������u̃}� u0��?���    j jEh@�h�h��� :�����   �  j$h�   �UR��(����3��} ���E܃}� uh�j jHh@�j�(������u̃}� u0�|?���    j jHh@�h�h��9�����   �  �U�U؋E؃x |�M؃9 s�3?���    �   ��  �U�UԋEԃx|"�Mԁ9�o@�v�?���    �   �  �&��j jRh@�h�h���U�R�-����P�%2����j jSh@�h�hx��E�P�;%����P��1����j jTh@�h�h<��M�Q�'/����P��1�����U�UЋEЃx ��   �MЁ9�� ��   �E���M�1+��Au�E�M�Q�UR�8�����E�}� t�E���  �}� tO�EP�#&������t?�E���M�+ȋE�M�E�M�Q�UR�7�����E�}� t�E��  �E�@    �  �MQ�UR�7�����E�}� t�E��`  �}� t7�EP�%������t'�M���ȋ�E�E��+��M�u�U�B    ��E� ��ȋ�E��+��M�u�j j<�U�R�E�P��%���M��U�: }�E���<�U�
�E��<�M�� �E�M�U�B�����j j<�E�P�M�Q��%�����u�}�j j<�U�R�E�P�u%���M�A�U�z }!�E�H��<�U�J�E��<�M�� �E�M�U�B�����j j<�E�P�M�Q�o%�����u�}�j j�U�R�E�P�%���M�A�U�z }!�E�H���U�J�E���M�� �E�M�j j�U�R�E�P�%���E�U�}� |D�}� v<�M�U�B���   ���E�P�M�UJ�E�H�M�UJ�E�H�   �}� ��   |
�}� ��   �M�Q�E�D��   ���E�P�M�U�B��E̋M�ỦQ�}� @�E�H���U�J�E�M�Q��m  �M�A�U�B   �E�H���U�J��E�MA�U�B3�_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����*���E��}� u3�� �EP�M�Q�4�����E��}� t3���E���]������������������̋�U����E�P�|�M��� �>ՋU���ޱ�j h��� RQ�8���E��U�}�|	�}��o@�v�E������E������} t�E�M���U�P�E��U��]�������������������������������������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uht�j jphP�j�.!������u̃}� u.�8���    j jphP�h0�ht��2��������)  �} t�} u	�E�    ��E�   �M̉MЃ}� uh�j jshP�j� ������u̃}� u.�8���    j jshP�h0�h�� 2��������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R��,�����E��} u�E��P�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj ��1�����EċE���]�������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP��3����]���������������̋�U��Q�M��EP�M�Q�f(������]� ����������������̋�U��Q�M��E�� ̤�M�Q�� ������]��������������̋�U��Q�M��M������E��t�M�Q�* �����E���]� �����������������̋�U��Q�M��EP�M�Q�f#������]� ����������������̋�U��Q�M��E�P�J1������]�������̋�U��Q�M��E���	P�M��	Q�]!�����������]� �������������������̋�U��Q�M��E���	P�M��	Q�!��������؋�]� ��������������������̋�U��Q�M��E���	P�M��	Q�� ����3҅���]� �����������������̋�U��Q�M��E�����]�������������̋�U��Q�M��E�� ̤�E���]� ��������������������̋�U��Q�M��E���]� ��������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̋�U����]����̋�U��Q�= 	 u� 	   ��= 	}
� 	   h�   hԤjj� 	P�2��������=�� u?� 	   h�   hԤjj� 	Q��1��������=�� u
�   �   �E�    �	�U����U��}�}�E������M���������E�    �	�E����E��}�}f�M����U����������<�t8�M����U����������<�t�M����U����������< u�M���ǁ�������3���]������������������������������������������������������������������������������������̋�U���������t���j���Q�!(����]�������������������̋�U��}��r4�}0�w+�E-������P�������M�Q�� �  �E�P��M�� Q��]�������������������������������̋�U��}}#�E��P�l�����M�Q�� �  �E�P��M�� Q��]�������������������̋�U��}��r4�}0�w+�E�H������U�J�E-������P�{&������M�� Q��]�������������������������������̋�U��}}#�E�H������U�J�E��P�&������M�� Q��]�������������������̋�U��E���]�����������������̋�U��Q����E��M�Q�l�E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�)����]����������������������̋�U��jh �j��+����h ���P��]����������������������̋�U���8  ���3ŉE��}�t�EP�p����ǅ����    jLj ������Q�������������U��� ����E��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �M�������U�������E�H��������U�������E�������M�������X�E�j ���U�R������������ u�}� u�}�t�EP�V�����M�3�������]�������������������������������������������������������������������������������������������������̋�U��Q�E�    ����E��M�Q�l�E��UR���E�E����E���]������������������̋�U��Q�E�    ����E��M�Q�l�E��E���]�����������������������̋�U��EP�MQ�UR�EP�MQ��&����]�������������̋�U��EP�MQ�UR�EP�MQ�(&��]����������������̋�U��V����M��UR���������3,���0^]������������������������̋�U��Q�E�    �	�E����E��}�-s�M��U;���u�E������7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]��������������������������������������������̋�U��Q�x���E��}� u	�   ���T+���M�3���]�������������������̋�U��Q3��} ���E��}� u!h��j h�   h(�j�������u̃}� u%j h�   h(�h�h���%�����   ���*���U� �3���]������������������������������������������̋�U��Q����E��}� u	�   ���+���M�3���]�������������������̋�U��Q3��} ���E��}� u!h��j h�   h(�j�������u̃}� u%j h�   h(�h��h���%$�����   �����U� �3���]������������������������������������������̋�U��Q����E��}� u	�8����E�����]���������̋�U��Q����E��}� u	�<����E�����]���������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uhЧj jahX�j�r������u̃}� u.��(���    j jahX�h$�hЧ��"��������h  3҃} �U؃}� uh��j jbhX�j�������u̃}� u.�o(���    j jbhX�h$�h���z"��������  j�������E�    �(��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�(�j�U�R�Y�����43�uh��j jhX�j�������u��E������c'���    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;(�tM�U�z t�E�H�U���M��E�H�J�U��    �E�(��H�(��E��M�(��h�   hL�jj�B	�����E�}� u�E������&���    �L�U��    �E�(��H�=(� t�(��E��M��A   �E�   �U�E�B�M�(��E������   �j�{����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP������E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR�\����]���������̋�U��X"  �^�����3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj ����u8j h<  hX�h�h��hT�h  ������R�*%����P������������E��M�Q�w������@v`�U�R�f�����M��TA��U�j hE  hX�h�hH�j���P�M�������+����  +���P�M�Q�l����P�<�����} t'�UR� ������@v�EP�������M�TA��U��#��� �������#���     �}uǅ����0��
ǅ����,��M���t�E�������
ǅ����,��M���t�}uǅ������
ǅ����,��E���tǅ������
ǅ����,��} t�U�������
ǅ����,��} tǅ������
ǅ����,��} t�E�������
ǅ����,��} tǅ����ܪ�
ǅ����,��}� t�M��������'�} t�U�������
ǅ����,��������������}� tǅ������
ǅ����,��} tǅ����Ī�
ǅ����,�������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M��<�Rh��h�  h   ������P�����D�E�}� }*j h`  hX�h�hةj"j�!���Q������ �!����������}� }8j hc  hX�h�h �h��h   ������P�"����P�����h  h`�������Q������������������uj�4����j���������u�   �3��M�3��!����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP�m���E]������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�������E��E�    �E���]�����������������̋�U���0�E� �E�   �E���E��M����M�U��B3���EԋM�Q�U�R��  ���E�H��f�   �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M��	���E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=�~ t h�~�#������tj�UR��~���M����U�����E��H;M�th���U�R�M����U��'���E��M�H�U�R�E�P��   ���U�M�I� �������&�U��z�th���E�P�M�������������E��M߅�t�U�R�E�P�   ���E��]������������������������������������������������������������������������������������������������������������������������̋�U����E�8�t%�M��E��M��U�EB3E��E��M�� ���M�Q�E��M��U�EB3E��E��M��������]���������������������������������̋�U��Q�EP�MQ�UR���P�MQ�������E��E���]������������������̋�U��j j j�EP�MQ�����]�������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�D   ���E��}� u�}� t������t
�����M���E���]������������������������̋�U��Q�EP�MQ�UR�EP�MQ�   ���E��}� t�E��?�} u�} t	�U�   �E��%�EP��������u�} t	�M�   3��뗋�]�����������������������������̋�U��j j j�EP������]�������̋�U��j�hȡh9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�l�����E�    �=�� vU�����9��u6������u!h��j h  hH�j�������u����    �������������E؃=���t�M�;��u̃=�� tu�UR�EP�M�Q�UR�EPj j�������uP�} t%�MQ�URh�j j j j �������u�� h�h�j j j j ��������u��D  �U����  ��t�����u�E�   �}�v3�MQh��j j j j�������u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t hx�h�j j j j�K������u̋M��$�MԋU�R��������E܃}� u�} t	�E�    �r  ���������}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+��;Mv���U����
����������E������;��v�������=�� t����M܉H�	�U܉���E܋����U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉��j���R�E܃�P�� ����j���Q�U�E܍L Q� �����UR���P�M܃� Q� �����U܃� �U��E������   �j�����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�(������E��}� u�}� t�����t
����U���E���]����������������������������̋�U��Q�} v�����3��u;Es�����    3��K�E�E�E�MQ�UR�EP�MQ���R�EP��������E��}� t�MQj �U�R�������E���]���������������������������������������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�l������E��}� u�}� t�����t
�����M���E���]������������������������̋�U��Qj j j�EP�MQ�UR��������E��E���]����������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    j�
������E�    j�EP�MQ�UR�EP�MQ�b   ���E��E������   �j�O
����ËE�M�d�    Y_^[��]����������������������������������������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R�������  �} t�}� u�EP�MQ�F
����3��  �=�� vV�����9��u6�������u!h��j h�  hH�j���������u����    �������������U�=���t�E�;��u̃=�� ty�MQ�UR�E�P�MQ�U�R�EPj�������uR�} t%�MQ�URh\�j j j j ���������u�� h0�h�j j j j ��������u�3��  �}��v`�} t)�UR�EP�M�Qh�j j j j�v����� ��u���E�Ph��j j j j�U�������u��!���    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh��j j j j���������u�� hx�h�j j j j���������u��Qj���R�E�����P�  ����t1�MQh �j j j j��������u��b���    3��t  �EP��������u!hȱj h  hH�j��������u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!h �j h#  hH�j�c�������u��d�M�Q����  ��u�E%��  ��u�E   �M���;Qs1�EPh�j j j j��������u��v���    3��  �} t%�U���$R�E�P�������E��}� u3��_  �#�M���$Q�U�R�������E��}� u3��:  3�u����������}� u|�=���s9�U���+B������+��;M�v���U�����
��������E����+H������U�������;��v�������U��� �U�E��M�;Hv$�U��E�+BP���Q�U��E�BP�h�����j���Q�U�U�R�O������}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!hh�j h�  hH�j�j�������u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8���;M�t!h,�j h�  hH�j��������u̋E��H����U��z t�E��H�U����7���;M�t!h�j h�  hH�j���������u̋E������=�� t����E��B�	�M�����U�����M��A    �U�����E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es����    3��g�E�E�E��} t�MQ�-������E��UR�EP�MQ�U�R�EP������E�}� t �M�;M�s�U�+U�Rj �E�E�P��������E��]����������������������������������������������������̋�U��Qj j j�EP�MQ�������E��E���]����������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    3��} ���E��}� u!h��j h�  hH�j�u�������u̃}� u-��
���    j h�  hH�h��h��������3��c�}�v�
���    3��Nj�?������E�    j �UR�EP�MQ�UR�EP�������E��E������   �j� ����ËE�M�d�    Y_^[��]�������������������������������������������������������������������̋�U��j�EP������]�����������̋�U��j�h(�h9�d�    P��SVW���1E�3�P�E�d�    j�J������E�    �EP�MQ�Y������E������   �j������ËM�d�    Y_^[��]����������������������������������̋�U��Q�=�� vU�����9��u6������u!h��j h  hH�j��������u����    ����������} u�l  �}uOj���P�M�����Q�	  ����t/�URh��j j j j��������u��}���    �  �=�� tDj j j �MQj �URj�������u%hp�h�j j j j �Y�������u���  �MQ�}�������u!hȱj h*  hH�j��������u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!h�j h0  hH�j�*�������u̋�����m  j���P�M���Q�k  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��`�Ph@�j j j j�A�����(��u��<�U��� R�E��HQ�U��B%��  ��`�Qh��j j j j������ ��u�j���P�M��Q�E��L Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��`�Phеj j j j������(��u��<�U��� R�E��HQ�U��B%��  ��`�Qh0�j j j j�I����� ��u̋E��xue�M��y����u	�U��z t!h��j hi  hH�j�o�������u̋M��Q��$R���P�M�Q��������U�R�Z������Q  �E��xu�}u�E   �M��Q;Ut!hP�j hw  hH�j���������u̋M����+Q����������   �M��9 t�U���M��Q�P�6���;E�t!h�j h�  hH�j��������u̋U��B����M��y t�U��B�M����5���;E�t!h�j h�  hH�j�M�������u̋U������M��Q��$R���P�M�Q�������U�R�.������(�E��@    �M��QR���P�M��� Q�u�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�EP�(�����]�����������̋�U��j�hH�h9�d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� u!h��j h�  hH�j�%�������u̃}� u1����    j h�  hH�h�h������������8  �=�� vV�����9��u6������u!h��j h�  hH�j��������u����    ���������j�������E�    �UR�B�������u!hȱj h�  hH�j�M�������u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!h�j h�  hH�j���������u̋E��xu�}u�E   �M��Q�U��E������   �j�[�����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������̋�U��Q����E��M����E���]������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    j��������E�    �EP�{�������te�M�� �M�U�B%��  ��tC�M�yt:�U�B%��  ��t*�M�yt!h�j h?  hH�j�K�������u̋E�M�H�E������   �j�������ËM�d�    Y_^[��]�������������������������������������������������������������̋�U��Q����E��M����E���]������������������̋�U�졜�]����̋�U��E�M���M��t�U�E��E���E;�t3���Ӹ   ]�����������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �����u
�   ��  j�������E�    �����E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$�x�h��h�j j j j �/�������u��   h��h�j j j j �
�������u��dhX�h�j j j j ���������u��Bh0�h�j j j j ���������u�� h��h�j j j j ��������u��E�    ��  �E�   ����E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��`��U���E��j���P�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh@�j j j j ������(��u��-�E�� P�M�QR�E�Ph��j j j j ������ ��u��E�    j���R�E�H�U�D
 P�2�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Phеj j j j ������(��u��-�U�� R�E�HQ�U�Rh0�j j j j ������� ��u��E�    �M�y ��   �U�BP���Q�U�� R��������ud�E�x t2�M�QR�E�HQ�U�� Rh0�j j j j �~����� ��u��"�M�� Qh��j j j j �Z�������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�Rh8�j j j j �	�����(��u��-�M�QR�E�� P�M�Qh�j j j j ������� ��u��E�    �G����E������   �j������ËE܋M�d�    Y_^[��]ÍI /���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    ����E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!h �j hy  hH�j�O�������u̃}� u0�����    j hy  hH�hػh �����������sj�+������E�    ����M�}�t7�U��t���   ��E��%��  ������    �M����E������   �j�K�����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������̋�U��j�hȢh9�d�    P���SVW���1E�3�P�E�d�    3��} ���E��}� u!h�j h�  hH�j���������u̃}� u+�6����    j h�  hH�h̽h��>������s�����u�fj�������E�    ����E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j�������ËM�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��3��} ��]����������������̋�U��} u3��1j j �E�� P��������u3���M�� Qj �l�R��]������������������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP��������u3���   j��������E�    �M�� �M��U��B%��  ��t"�M��yt�U��B%��  ��t	�M��yukj�UR�EP�o�������tU�M��Q;UuJ�E��H;��<�} t�U�E��H�
�} t�U�E��H�
�} t�U�E��H�
�E�   ��E�    �E������   �j������ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U��Q�EP�8�������u�����M�� �M��U��B��]������������������̋�U��Q����E��M����E���]������������������̋�U����]����̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� u!hȾj h�  hH�j��������u̃}� u.������    j h�  hH�h��hȾ��������m  j�s������E�    �U�����E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡ���E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�RhP�j j j j ������� ��u���M�Qh(�j j j j ���������u������E����H,�U����B0�E������   �j������ËM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���V�E�    3��} ���E�}� u!hȾj h�  hH�j��������u̃}� u0�x����    j h�  hH�h<�hȾ������3��  3҃} �U��}� u!h�j h�  hH�j��������u̃}� u0�����    j h�  hH�h<�h�������3��0  3Ƀ} ���M�}� u!h�j h�  hH�j�E�������u̃}� u0�����    j h�  hH�h<�h�������3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u�����t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M��x����M�����P�MQ�#   ���M��z�����]��������������������̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    �E�    j�C������E�    h`�h�j j j j ��������u̃} t�M��U����E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u�����u��  �U�z twj j�E�HQ�v�������tj�U�BP����t$�M�QRhH�j j j j ���������u��)�M�QR�E�HQh8�j j j j ��������u̋E�HQh0�j j j j ��������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph�j j j j �6����� ��u̃=�� t,j�U�� R����u�E�HQ�U�� R�������E�P�MQ�  ���   �U�zu;�E�HQ�U�� Rh��j j j j ��������u̋M�Q�UR�x  ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� Ph��j j j j �^����� ��u̋U�R�EP�  ��������E������   �j�7������hh�h�j j j j ��������u̋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���t���3ŉE��EP�M��U����E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M�������t3�M���������   ~ �M��{���PhW  �E�P��������E��hW  �M�Q�M��Q���P�������E��}� t	�U��U���E�    �E��M��L��!�����U������     �E�Ph���M�k��1   +�R�E�k��L�Q���������}*j h	  hH�h��hةj"j������R������ �����M��������U��D� �E�P�M�Qhx�j j j j ��������u̍M������M�3�������]������������������������������������������������������������������������������������������������������������������̋�U���8���3ŉE��E�P�%������}� u�}� u�����t7�}� t1h��h�j j j j ���������u�j �S������   �3��M�3�������]������������������������������������̋�U���3��} ���E��}� u!hȾj h�	  hH�j��������u̃}� u.�����    j h�	  hH�hT�hȾ�������   �E�    �	�U����U��}�}>�E���`�Q�U��E�L�Q�U��E�L�Qh0�j j j j ������� ��u�볋E�H,Qh�j j j j ��������u̋E�H0Qh��j j j j �|�������u̋�]�������������������������������������������������������������������̋�U��j j j �EP�MQ�_�����]�������������������̋�U��EP�MQj �UR�EP�+�����]���������������̋�U��j j j �EP�MQ�UR������]���������������̋�U��j j j �EP�MQ�UR�EP������]�����������̋�U��EP�MQj �UR�EP�MQ�Q�����]�����������̋�U��EP�MQj �UR�EP�MQ�UR������]�����������������������̋�U��j j �EP�MQ�UR�-�����]�����������������̋�U���(�E��#E������E�u!h�j h�
  hH�j���������u̃}� u0�]����    j h�
  hH�h��h��e�����3��@  �} t�U;Ur	�E�    ��E�   �E܉E��}� u!h��j h�
  hH�j�{�������u̃}� u0������    j h�
  hH�h��h���������3��   �}v�U�U���E�   �E؃��E3�+M���M�U�E�L�M��UU��U�E;E�v�e����    3��i�MQ�URj�E�P��������E�}� u3��F�M�M�M�U��#�+M�M��E�+E���E�j���Q�U���R�������E��M��E���]������������������������������������������������������������������������������������������������������������������������̋�U��j j �EP�MQ�UR�EP������]�������������̋�U��j j �EP�MQ�UR�EP�MQ�������]���������̋�U���4�} u!�EP�MQ�UR�EP�MQ�`������  �} u�UR�P�����3��  �E������E�j���Q�U��R��������t1�EPh��j j j j��������u������    3��C  j���R�E���P�X�������u�MQh��j j j j�g�������u̋E��#E������E�u!h�j h�  hH�j��������u̃}� u0������    j h�  hH�h<�h��������3��  �} t�U;Ur	�E�    ��E�   �EԉE؃}� u!h��j h�  hH�j��������u̃}� u0�v����    j h�  hH�h<�h���~�����3��  �U��P�q������M��U++E�}v�E�E���E�   �MЃ��M3�+U���U�E�M�T�U�EE�E�M;M�v������    3��   �UR�EPj�M�Q�<������E��}� u3��   �U�U�U�E��#�+U�U��M�+M���M�j���R�E���P�������M��U���E�;Ev�M�M���U�ŰE�P�MQ�U�R�2�����j�E��Q��������E���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�    �E�    �} v�����3��u;Es�/����    3��s�E�E�E��} t�MQ�UR�EP�w������E��M Q�UR�EP�MQ�U�R�EP�������E�}� t �M�;M�s�U�+U�Rj �E�E�P��������E��]��������������������������������������������������������̋�U��EP�������]�������������̋�U��Q�} u�   �E������E�j���Q�U��R��������t!�EPh �j j j j�,�������u��Lj���R�E���P���������u�MQh��j j j j���������u�j�E��Q�u�������]�����������������������������������������������������̋�U��Q����E��M����E���]������������������̋�U��Q����E��E���]�����������̋�U����]����̋�U��EP�MQ�UR�������]���������������������̋�U��� �E�    �E�    �E�    �E�    �E�    3��} ���E�}� u!h��j h�  hH�j��������u̃}� u.�}����    j h�  hH�ht�h������������w�E�    �U������U��E��Q�g������E��U��E+�E�3�+M���M�}v�U�U���E�   �E����E�M�U�D
+E�E�M�+M�+M�M��E���]�������������������������������������������������������������������̋�U��j�hH�h9�d�    P���SVW���1E�3�P�E�d�    �}�u�����     �N���� 	   ����  �} |�E;h�s	�E�   ��E�    �M؉M��}� uh8�j j.h��j��������u̃}� u9�����     ������ 	   j j.h��h��h8������������  �E���M���������D
������؉E�uh��j j/h��j��������u̃}� u9�����     �Y���� 	   j j/h��h��h���d���������   �UR�������E�    �E���M���������D
��t�MQ�������E��4������ 	   �E�����3�uh��j j9h��j�L�������u��E������   ��MQ菽����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QV�EP�q��������t]�}u������   ��u�}u(����HD��tj�6�������j�*�����;�t�UR������P����t	�E�    �	���E��EP�(������M���U���������D �}� t�M�Q����������3�^��]����������������������������������������������������̋�U��Q3��} ���E��}� uh�j j)h��j�T�������u̃}� u+�����    j j)h��h��h�������������U�B��]�������������������������������̋�U��} uh��j j.h8�j�Ѿ������u̋M�Q��   tK�E�H��t@j�U�BP��������M�Q�������E�P�M�    �U�B    �E�@    ]��������������������������������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    �} uj �  ���@�EP�C������E�    �MQ�H������E��E������   ��UR�6�����ËE�M�d�    Y_^[��]������������������������������������������̋�U��} uj �n  ���@�EP��������t����+�M�Q�� @  t�EP�X�����P����������3�]�����������������������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R�������P�P�����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����������������������������������������������������̋�U��j�   ��]���������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�ܼ�����E�    �E�    �	�E����E��M�; 	��   �U����<� ��   �M�������H��   ��   �U�����Q�U�R�������E�   �E�������B%�   te�}u%�M������P�|��������t	�M���M��:�} u4�U������Q��t!�E������R�>��������u�E������E�    �   ��E������R�E�P��������������E������   �j�-�����Ã}u�E����E܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������̋�U���V�E�    3��} ���E��}� uh`�j jih��j躹������u̃}� u.�����    j jih��h��h`��&����������  �U�U��E��H��   t�U��B��@t����  �M��Q��t�E��H�� �U��J����  �E��H���U��J�E��H��  u�U�R��������E��M��Q��E��HQ�U��BP�M�Q������P�&������U��B�E��x t	�M��y�u.�U��B��������M�A�U��B�E��@    �����   �M��Q��   u�E�P���������t@�M�Q���������t/�U�R�v����������E�P�e�������������E���E����M��Q��   ���   u�E��H��    �U��J�E��x   u#�M��Q��t�E��H��   u
�U��B   �E��H���U��J�E������   �U��E�����U��
�E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������̋�U���p�E�P��h�   h|�jj@j �������E��}� u�����  �M�����h�    �	�U���@�U����   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E����  �}� ��  �M��U��E���E��M�M��M��}�   }�U��U���E�   �E��E��E�   �	�M����M��h�;U���   h�   h|�jj@j �o������E��}� u�h��E��   �M��U������h��� �h��	�M���@�M��U�����   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tv�U����u�M��R����t[�E����M���������M��U��E���
�U��E���Jh�  �U���R����u����`  �E��H���U��J�;����E�    �	�E����E��}��!  �M������M��U��:�t�E��8���   �M��A��}� u	�E�������U�����҃���U��E�P���E��}����   �}� ��   �M�Q���E��}� tr�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P����u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A������h�R��3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �	�E����E��}�@}y�M��<��� tg�U������E��	�M���@�M��U�����   9E�s�M��y t�U���R����j�E�����Q覿�����U�����    �x�����]���������������������������������������������������̋�U���T�t��E��E�    �E�    �E�    �} uh �j jDh��j��������u̃} uhp�j jEh��j轰������u̃} uh`�j jFh��j虰������u̋M��� u�E���E��M��UĀ}�at8�}�rt�}�wt�<�E�    �E���E��   �E�  �M���M��   �E�	  �U���U��q3�t	�E�   ��E�    �M��M܃}� uh(�j jbh��j��������u̃}� u-�N����    j jbh��h�h(��Y�����3��  �E�   �E���E�M����7  �}� �-  �E��M��U��� �U��}�T��  �E�����$����  �U��t	�E�    �'�E���E�M����M�U�ʀ   �U�E����E��  �M�� �  t	�E�    ��U�� �  �U��  �E�% �  t	�E�    ��M�� @  �M��p  �}� t	�E�    ��E�   �U�� @  �U��I  �}� t	�E�    ��E�   �E�%�����E��#  �}� t	�E�    ��E�   �M�� �M���   �}� t	�E�    ��E�   �U���U���   �E�%   t	�E�    ��M��   �M��   �U��@t	�E�    �	�E��@�E��   �M�ɀ   �M��   �E�   �E�    �w3�t	�E�   ��E�    �E��E؃}� u!h(�j h�   h��j蠭������u̃}� u0�����    j h�   h��h�h(��	�����3��i  �����}� �h  �U��� u�M���M��j�URh����������tw3�t	�E�   ��E�    �M��Mԃ}� u!h(�j h�   h��j��������u̃}� u0�N����    j h�   h��h�h(��V�����3��  �E���E�M��� u�E���E��M���=tw3�t	�E�   ��E�    �M��MЃ}� u!h(�j h�   h��j�L�������u̃}� u0�����    j h�   h��h�h(�赽����3��  �E���E�M��� u�E���E��jh���MQ�è������u�U���U�E�   �E���   jh���MQ蓨������u�U���U�E�   �E��   jh���MQ�c�������u�U���U�E�   �E��w3�t	�E�   ��E�    �U��Ũ}� u!h(�j h  h��j�)�������u̃}� u0�����    j h  h��h�h(�蒼����3���   �M��� u�E���E��M���҃��U�u!h��j h  h��j說������u̃}� u-�����    j h  h��h�h��������3��vh�  �MQ�U�R�EP�M�Q�`�������t3��Q���������E�E��M��U�Q�E��@    �M��    �U��B    �E��@    �M��U��Q�E���]ÍI �Yx�5W��|� 	
����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E�    j�S������E�    �E�    �	�E���E�M�; 	�z  �U����<� ��   �M������H��   ��   �U������Q�� �  ��   �}�~�}�}�E��P荢������u�  �M�����P�M�Q�п�����U������Q��   t�E�����R�E�P臶�����0����M������E��   �   jYh(�jj8�������E܋M����E܉��}� twh�  �M������� P����u)j�M�����P�������M�����    �6�E������� R���E������U��E��@    ��n����}� tC�M��Q�� �  �E��P�M��A    �U��B    �E��     �M��A    �U��B�����E������   �j�ղ����ËE��M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������SVW�T$�D$�L$URPQQh�#d�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�t����   �C賥���d�    ��_^[ËL$�A   �   t3�D$�H3��l���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�Ѵ��3�3�3�3�3���U��SVWj Rh6$Q耮��_^[]�U�l$RQ�t$������]� ���������������������������������������������������������������������������������������������̋�U����} uh`�j j?h��j螢������u̋M�M��U�R蠫����P�ϴ������u3��  ������� 9E�u	�E�    �������@9E�u	�E�   �3���   ���������M��Q��  t3��   �E��<�� u\j[hd�jh   �������E�M��U����}� u0�E����E��M��U��Q�E��M���U��B   �E��@   �/�M��U�����A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]��������������������������������������������������������������������������������������̋�U��Q�} t'�}t!h�j h�   h��j��������u̋M�M��} tG�U��B%   t:�M�Q�������U��B%�����M��A�U��B    �E��     �M��A    ��]��������������������������������������̋�U���   ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M������E�    �u����E�3Ƀ} �������������� u!h�j h  h��j�͟������u̃����� uF�+����    j h  h��h��h��3�����ǅ ��������M�職���� �����  �E�������������Q��@��   ������P�h������������������t-�������t$���������������������������
ǅ�����������H$�����х�uV�������t-�������t$���������������������������
ǅ�����������B$�� ���ȅ�tǅ ���    �
ǅ ���   �� ��������������� u!h`�j h  h��j�X�������u̃����� uF趵���    j h  h��h��h`�辯����ǅ��������M�����������U  3Ƀ} �������������� u!ht�j h  h��j�Н������u̃����� uF�.����    j h  h��h��ht��6�����ǅ��������M�脵���������  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���g  ������ �Z  �������� |%��������x��������H����������
ǅ����    ���������������������������h�����������������������������  �������$��8�E�    �M������P������R�ǝ��������   ������P�MQ������R�t  ���E��������U���U����������؉�����u!hh�j h�  h��j��������u̃����� uF�o����    j h�  h��h��hh��w�����ǅ��������M��ų��������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK��������9�$��8�E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP�������E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ辯�����Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  ��������49�$� 9�E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ���������9�$�d9�U���0  u�E�   �E��M���  tUǅ|���    �UR腨����f������������Ph   ������Q�U�R��������|�����|��� t�E�   �&�EP虭����f��x�����x����������E�   �������U��W  �EP�e�������t�����t��� t��t����y u� ��U��E�P�������E��P�M���   t&��t����B�E���t�����+����E��E�   ��E�    ��t����B�E���t�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������l����MQ蒬�����E��U���  te�}� u���E��E�   �M���h�����l�����l�������l�����t��h������t��h�������h����ɋ�h���+M����M��[�}� u	� ��U��E���p�����l�����l�������l�����t��p������t��p�������p����ɋ�p���+E��E��  �MQ賫������d����Ѣ������   3�tǅ����   �
ǅ����    ��������`�����`��� u!h�j h�  h��j��������u̃�`��� uF�y����    j h�  h��h��h�聧����ǅ��������M��ϭ��������  ��  �U��� t��d���f������f����d�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  h��j�Ú�]  R�������E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���X�����\����M��#���P�E�P�M�Q������R�E�P�M�Q��X���R�H�P�l�Ѓ��M���   t$�}� u�M��ٓ��P�U�R�T�P�l�Ѓ���������gu*�U���   u�M�褓��P�E�P�P�Q�l�Ѓ��U����-u�M���   �M��U����U��E�P�������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ蠙������H�����L����   �U���   t�EP�x�������H�����L����   �M��� tB�U���@t�EP�7���������H�����L�����MQ�����������H�����L����=�U���@t�EP����������H�����L�����MQ�ڧ����3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��M̋Ũ��U̅���@����D���t{�E��RP��D���Q��@���R������0��T����E��RP��D���P��@���Q蒧����@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �J  ���U�R������P�MQ�U�R�E�P�{  ���M���t$�U���u������P�MQ��<���Rj0��  ���}� ��   �}� ��   ǅ$���    �E���8����M܉�4�����4�����4�������4�������   ��8���f�f������������Pj��(���Q��0���R��������$�����8�������8�����$��� u	��0��� uǅ���������*�M�Q������R�EP��0���Q��(���R�z  ���V�����E�P������Q�UR�E�P�M�Q�T  �������� |$�U���t������P�MQ��<���Rj ��  ���}� tj�E�P�������E�    �v���������������M�貦��������M�3��L�����]��*�+,�,�,�,-W.Z,e,O,D,r,{, �I �-<.Y-G.R. ��1�.�/�3>/�1�.�3�0�3�3�/�3�3�6   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�Z������E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A�]��������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U��E����U�
�E�f�A�]�������������������̋�U��j�hأh9�d�    P���SVW���1E�3�P�E�d�    詒���� �E�3��} ���E؃}� uht�j j4h@�j��������u̃}� u+�N����    j j4h@�h�ht��Y���������i�U�R��������E�    �E�P�.������E܋MQ�UR�EP�M�Q�U���E��U�R�E�P�`������E������   ��M�Q�Õ����ËE��M�d�    Y_^[��]�����������������������������������������������������������������������̋�U��EP�MQ�URh(�覂����]����������������̋�U��EP�MQ�URh:��v�����]����������������̋�U��EP�MQ�URh��F�����]����������������̋�U��EPj �MQh(�������]������������������̋�U��EPj �MQh:�������]������������������̋�U��EPj �MQh�踁����]������������������̋�U���(  ���������5��=�f�0�f�$�f� �f���f�%��f�-����(��E ���E� ��E�,��������h�  � �����	 ���   �������������������X�`�j������j ��h�����=`� u
j������h	 ���P����]����������������������������������������������������������������������������������̋�U��j ��]�����������������̋�U����]� ����������������̋�U��EP��Q����]� �������������������̋�U���]����̋�U��Q��P���E��}� u ���Q�l�E��U�R��P���E���]������������������������������̋�U��EP�MQ���R�l��]� ���������������̋�U���h8����E��}� u�F���3���  h,��E�P�T���h��M�Q�T���h��U�R�T���h ��E�P�T����=�� t�=�� t�=�� t	�=�� u,�������������������������=��t���Q��R����u3���   耄�����P��������Q��������R��������P������T�����u����3��   h����Q�l�У��=��u	����3��rh  h��jh  j�k������E��}� t�U�R��P���Q�l�Ѕ�u	蛈��3��(j �U�R�?������h�M���U��B�����   ��]������������������������������������������������������������������������������������������������������������������������������������̋�U��=��t��P���Q�l���������=��t��R���������Ny��]����������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    h8����E�E�@\���M�A    �U�B   �E�@p   �MƁ�   C�UƂK  C�E�@h`�j������E�    �M�QhR���E������   �j�_������j��~�����E�   �E�M�Hl�U�zl u�E�D��Hl�U�BlP�z������E������   �j������ËM�d�    Y_^[��]��������������������������������������������������������������������������̋�U������E���P�Av���ЉE��}� u}j h�  h��jh  j�~�����E��}� tW�M�Q��R���P�l�Ѕ�t%j �M�Q�E������h�U���E��@�����j�M�Q蟊�����E�    �U�R���E���]�����������������������������������������������������������̋�U��Q�w���E��}� u
j�o������E���]�����������̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P��������M܃y, tj�U܋B,P覉�����M܃y4 tj�U܋B4P茉�����M܃y< tj�U܋B<P�r������M܃y@ tj�U܋B@P�X������M܃yD tj�U܋BDP�>������M܃yH tj�U܋BHP�$������M܁y\��tj�U܋B\P������j��{�����E�    �M܋Qh�U��}� t%�E�P����u�}�`�tj�M�Q������E������   �j�������j�{�����E�   �U܋Bl�E�}� t4�M�Q��������U�;D�t�}�@�t�E�8 u�M�Q�v�����E������   �j謇�����j�U�R�.������M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������̋�U��=��tO�} u)��P����t��Q��R���ЉEj ��P���Q�l�ЋUR莄���=��tj ��P��]������������������������������������������̋�U���h]���̋�U����]���̋�U��Q�=� th��ɋ������t�EP�����C���hwh�t�������E��}� t�E��Gh��lx����h�sh p�R  ���=d� thd��^�������tj jj �d�3���]���������������������������������������������������̋�U��j j �EP�>  ��]���������̋�U��j j�EP�  ��]���������̋�U��jj j �   ��]�����������̋�U��jjj ��  ��]�����������̋�U��蘉���EP�z����h�   �y��]��������������̋�U��Q� ��E��	�M����M��}� t�U��: tj�E��Q��������j� �R������� �    ����E��	�M����M��}� t�U��: tj�E��Q�Ǆ������j���R贄�������    j���P蚄����j���Q艄����j�\�R�lP�q��������    ���    ��{���\����P����u'�=��`�tj���Q�&��������`����R����]�����������������������������������������������������������������������������������������������̋�U��j�hX�h9�d�    P���SVW���1E�3�P�E�d�    �ڄ���E�    �=��U  ��   �E���} ��   �\�Q�l�E�}� ��   �X�R�l�E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r�Pz���U�9u��E�;E�s�h�M؋R�l�E��)z���M؉�U܋\�R�l�EСX�P�l�E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��T���h({hx�A  ��h0}h,|�/  ���=� u#j��us������ t��   �m���Ā���E������   ��} t�^n��Ã} t���   �Fn���MQ�bv�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������̋�U���hl����E��}� thX��E�P�T�E��}� t�MQ�U���]�����������������̋�U��EP�n�����MQ��]�������������������̋�U��j�s����]���������������̋�U��j������]���������������̋�U��Q��w���E��E�P�4������M�Q�^������U�R�{�����E�P�k�����M�Q�ut�����U�R�z������]����������������������̋�U��E;Es�M�9 t�U��ЋM���M��]�����������������������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�����������������̋�U���3��} ���E��}� u!h��j h�  h��j�q������u̃}� u0�p����    j h�  h��h��h���x������   �y3҃=� �U��}� u!h��j h�  h��j�p������u̃}� u0�����    j h�  h��h��h���������   ��M���3���]������������������������������������������������������������������̋�U���3��} ���E��}� u!h��j h�  h��j��o������u̃}� u0�@����    j h�  h��hp�h���H������   �y3҃=� �U��}� u!hH�j h�  h��j�so������u̃}� u0�Ԇ���    j h�  h��hp�hH��܀�����   ��M���3���]������������������������������������������������������������������̋�U����=`� u��i���E�    ����E��}� u����e  �M����t,�E����=t	�U����U��E�P�q�����M��T�U���juh`�jj�E���P�	������E�M����=�� u�����   ����U��	�E�E��E��M������   �E�P�'q�������E��M����=��   j~h`�jj�E�P蒄�����M��U�: uj���P�|�������    ����rj h�   h��h��h���M�Q�U�R�E�Q������P�[x�����U���U��B���j���P�{�������    �M��    �H�   3���]��������������������������������������������������������������������������������������������������������������������̋�U����E�    �=`� u��g���4� h  h0�j �Ph0��h�����=	 t�	���t�	�U���E�0��E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   h��j�M��U���P��e�����E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�   ���U�������E����3���]�������������������������������������������������������������������������̋�U��E��]�����������������̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q�x������t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P�0v������t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R��u������t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    ���E��}� u3���   �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j ���E��}� tjJh��j�M�Q�h`�����E�}� u�U�R��3��Dj j �E�P�M�Q�U�R�E�Pj j ����uj�M�Q�lt�����E�    �U�R���E��]������������������������������������������������������������������������̋�V�؜��=؝s���t�Ѓ���؝r�^����������̋�V�����=��s���t�Ѓ�����r�^����������̋�U��Q�E�   j h   j � �l��=l� u3���   ��]�������������������������̋�U��l�P��l�    ]�������������������̋�U��=l� uh��j jhh�j��d������u̡l�]�������������̋�U����E�    �E�    �=��N�@�t���%  ��t����щ���   �U�R�|�E��E�M�3M��M��3E�E��h3E�E��3E�E�U�R��E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E�G  ��E�E�M����U��҉����]����������������������������������������������������������������̋�U��}csm�u�EP�MQ�&w������3�]����������̋�U�����^���E��}� u3���  �E��H\Q�UR�S  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����v  �E��H`�M�U��E�B`�M��y�4  �0��U��	�E����E��0�4�9M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]��������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��;Ut�E����E��<�k�M9M�s�ڋ<�k�U9U�s
�E��;Mt3���E���]������������������������̋�U��E��w$����������tRP�EQP�D   ��]ú`�R�   P�E�   QP�$   ��]�������������������������������̋�U���@  ���3ŉE��ES�]VW�}S������������ǅ����    ��\������������uS��w�����������5j j j�Wj h��  ��=   s&P������Qj�Wj h��  �օ�t�������������
ǅ������h  ��  ����������t%����������PSQW�}  �����"  2��������� ������u���  ��t�X����   h  ������R������Ph  ������Q���S�p������t-������������RWh��������P�EQ������RP���   �=�j j h
  ������Qj�������Rj h��  ����ׅ�t������j j h
  ������Pj�������Qj h��  �h��ׅ�t������������������������R�UPh@�VQSR����������u̋M�_^3�[�X����]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hx�h9�d�    P��$SVW���1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@��	�   Ëe��E������E�M�d�    Y_^[��]��������������������������������������̋�U��j�h��h9�d�    P��$SVW���1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@��	�   Ëe��E������E�M�d�    Y_^[��]����������������������������������������������������̋�U���  ���3ŉE��= ���E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ����������A��u�Њ@��u�W������+�O�OG��u��������ȃ�����Ȋ@��u�������+���O�OG��u������ȃ��_��l�� �������SjPQ�������^[�M�3��U����]��������������������������������������������������������������������̋�U���D  ���3ŉE�S�(�V�uW�}�����������   h��� ����   h��P�T�p�����   ����   �M�Vh��Qh����$Rh���~ Whx�h �������h�Q�ЋV��$RW�E�P�M�Q��   ��8h��U�Rh��E�Ph��������Q�������R�p�������������PjSQ������(_^[�M�3��?T����]�h��jSW�������M�_^3�[�T����]�����������������������������������������������������������������������������̋�U����ESV�u�E��EW3�+ƉE����M��r�   ;�s&�0�U���Qh��R�p��E��E����GF�ɋM�E�y� � _^[��]���������������������������������̋�U���  ���3ŉE��=$���E��   SV����   �ȍq�A��u�+΃�:��   ww������3Ɋ���������A��u�Њ@��u�W������+�O�OG��u��������ȃ�����Ȋ@��u�������+���O�OG��u������ȃ��_�����$�SjP�EP������^[�M�3��WR����]�����������������������������������������������������������������������̸   ����������̋�U��E��w	���]�3�]������̋�U��M��w�U������]Ã��]�����������̋�U��M�t��t��x�    ]�����������������̋�U��M�x��x��t�    ]�����������������̡t�����������̡x������������u�U��� PRSVWhp�hk�jBh �j��V������u�_^[ZX��]������������������������̋�U���]����̋�U��q�]�����f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U��������������������������������������������������������̋�U��j
�$�<�3�]����������̋�U��j jh(�h��hx�h   h   j �'e����P�_����]�������������������������̋�U��j �EP�$h����]�����������̋�U����EP�M��_^���M�R�Wd������et�E���E�M�R��S������u�E�Q�'d������xu	�U���U�E��M��M��S������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M���k����]������������������������������������������������̋�U��j �EP�'T����]�����������̋�U���V�EP�M��N]���M���t*�E�0�M���R������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��7R������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M��zj��^��]�������������������������������������������������������������������̋�U��Q�E�������Az	�E�   ��E�    �E���]���������������������̋�U����} t$�EP�MQ�U�R��T�����E�M���U��P��EP�MQ�U�R�[�����E�M���]������������������������������̋�U��j �EP�MQ�UR��g����]�������������������̋�U���D���3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�=c����3Ƀ} ���Mă}� u!hl�j h�  h��j��P������u̃}� u3�Gh���    j h�  h��h��hl��Ob�����   �  3�;E��ىM�u!h��j h�  h��j�~P������u̃}� u3��g���    j h�  h��h��h����a�����   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P�WI�����Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3��DJ����]��������������������������������������������������������������������������������������������������������������������̋�U���@�E�    �E P�M���X��3Ƀ} ���M܃}� u!hl�j h3  h��j��N������u̃}� u@�=f���    j h3  h��h��hl��E`�����E�   �M��f���E���  3�;E��ىM�u!h��j h4  h��j�gN������u̃}� u@��e���    j h4  h��h��h����_�����E�   �M��!f���E��}  3��} ����#E��	;E��ىM�u!hh�j h<  h��j��M������u̃}� u@�Ce��� "   j h<  h��h��hh��K_�����E�"   �M��e���E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�6  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��L������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h_  h��h��h��h���U�R�E�P�Be����P�W�����M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE�������t �U����0uj�M��Q�U�R�T�����E�    �M��c���Eċ�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�C����]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M���S���} }�E    3Ƀ} ���M��}� u!hl�j h�  h��j��I������u̃}� u@�9a���    j h�  h��ht�hl��A[�����E�   �M��a���E���  3�;E��ىM�u!h��j h�  h��j�cI������u̃}� u@��`���    j h�  h��ht�h����Z�����E�   �M��a���E��g  �E�  �M��;M��ډU�u!h�j h�  h��j��H������u̃}� u@�E`��� "   j h�  h��ht�h��MZ�����E�"   �M��`���E���  �M��Q�4�2`��%�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ��P�����E��}� t�U� �E��E��M��`���E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ�J�����E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M��~_���E���  �M��Q�?�_������ ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4�^��%�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M��E������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U��D���E�U��E܅���   �} ~}�M��Q���� #E�#U��M��V]��f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U��]���E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M���\��f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4��[��%�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�D������0�M��U���Uj h�  �E�P�M�Q�C���E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q�C���Ѓ�0�E��M���Mj jd�U�R�E�P�FC���E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�_C���ȃ�0�U�
�E���Ej j
�M�Q�U�R��B���E��U��E���0�M��U���U�E�  �E�    �M��Z���E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�9����]�����������̋�U���D���3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�mR����3Ƀ} ���Mă}� u!hl�j h*  h��j�@������u̃}� u3�wW���    j h*  h��h��hl��Q�����   ��   3�;E��ىM�u!h��j h+  h��j�?������u̃}� u3�W���    j h+  h��h��h���Q�����   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP�8�����Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�   ���EȋEȋM�3��9����]�����������������������������������������������������������������������������������������������������������̋�U���4�E�H���M��UR�M��3H��3��} ���E�}� u!hl�j h�  h��j�'>������u̃}� u@�U���    j h�  h��h��hl��O�����E�   �M���U���E��  3�;U��؉E�u!h��j h�  h��j�=������u̃}� u@�U���    j h�  h��h��h���O�����E�   �M��lU���E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P��  ���M��0�U����U���E�M�H�M��} ��   j�U�R�  ���M��'<��� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�  ���EPj0�M�Q��<�����E�    �M��%T���EЋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�R����]���������������̋�U���P���3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P�9M����3Ƀ} ���M��}� u!hl�j ho  h��j��:������u̃}� u3�CR���    j ho  h��h��hl��KL�����   �i  3�;E��ىM�u!h��j hp  h��j�z:������u̃}� u3��Q���    j hp  h��h��h����K�����   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R�Z3�����E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�_������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ��������M�3���3����]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�mP����]�����������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�K1�����E��{�}fu!�E P�MQ�UR�EP�MQ�LO�����E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ��0�����E��#�U R�EP�MQ�UR�EP�MQ�O�����E��E���]������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�UR�l1����]�����������������������̋�U��} t#�EP�.:������P�MQ�UUR��?����]����������������̋�U��Q�E�    �	�E����E��}�
s�M���0�R���M���0��ԋ�]������������������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y��������������������������������������������������������������������������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�j jh��j�5������u̃}� u0�mL���    j jh��h|�h��xF�����   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U�E�Ph�   �M��Q��4����3҃} �U��}� uhL�j jh��j�G4������u̃}� u0�K���    j jh��h|�hL��E�����   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q��3��������t3�t	�E�   ��E�    �M܉M�}� uh��j jh��j�,3������u̃}� u-�J��� "   j jh��h|�h���D�����"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9��s
����E���M+M����U+щU؋E�Ph�   �M+M��U�D
P�3����3���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    ��9���E��E��Hp#��t�U��zl ��   j�2�����E�    �E��Hh�M�U�;��tI�}� t%�E�P����u�}�`�tj�M�Q�W?�����Uࡈ��Bh����M�U�R���E������   �j�>������	�E��Hh�M�}� u
j �FD�����E�M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�hؤh9�d�    P���SVW���1E�3�P�E�d�    �E������8���E��[A���E܋Hh�M��UR��  ���E�E��M;H�  hN  h|�jh   ��)�����E��}� ��  �U܋rh��   �}��E��     �M�Q�UR�a1�����E؃}� ��  �E܋HhQ����u�U܁zh`�tj�E܋HhQ�=�����U܋E��Bh�M܋QhR���E܋Hp���-  ������  j�a0�����E�    �E��H����U��B����M��Q����E�    �	�E���E�}�}�M�U�E�f�TPf�M�����E�    �	�E���E�}�  }�M�M�U�A�������E�    �	�M���M�}�   }�U�U�E䊊  �����׋��R����u�=��`�tj���P�<�����M�����U�R���E������   �j��;������(�}��u"�}�`�tj�E�P�D<�����yE���    ��E�    �E؋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hX.d�    P��$���3�P�E�d�    �E�    �E�P�M���6���E�    ���    �}�u)���   �,�E��E������M��D���E��}�c�}�u)���   �(�E��E������M��D���E��N�4�}�u.���   �M���+����Q�U��E������M��ZD���E���E�E��E������M��@D���EЋM�d�    Y��]����������������������������������������������������������������������������̋�U���,���3ŉE�V�EP�������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0����;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E��� ��M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E������UU��B��MM��A����v����U�E�B�M�A   �U�BP��  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��p��f�DJ�ӋMQ�C  ��3��  �����} t!�}��  t�}��  t�UR�4��u����k  �E�P�MQ�0���9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�\  ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���=�� t�EP�  ��3�����^�M�3��K#����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���  �M��}�w-�U�����$���  ��  ��  �	�  �3���]ÍI ߟ������ ������������������������������������̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U���|��A���E�    �	�M����M��}�   }�UU��E���}���  �׋�]���������������������������������������������������������̋�U���(  ���3ŉE�������P�M�QR�0���-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj �o1���� j �M�QRh   ������Ph   ������Qh   �U�BPj �2����$j �M�QRh   ������Ph   ������Qh   �U�BPj ��1����$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�P�M���+���M��R!���H�y t �M��A!���P�B�E�M��9���E����E�    �M��9���E���M��9����]������������������������������������̋�U��=`� uj��:�����`�   3�]����������̋�U��Q�EP���M���    t�U���   P���M���    t�U���   P���M���    t�U���   P���M���    t�U���   P���E�    �	�M����M��}�m�U����E�|H��t$�M����U�|
P t�E����M�TPR���E����M�|L t$�U����E�|T t�M����U�D
TP��넋M���   �´   R����]���������������������������������������������������������������������������������̋�U��Q�} �  �EP���M���    t�U���   P���M���    t�U���   P���M���    t�U���   P���M���    t�U���   P���E�    �	�M����M��}�m�U����E�|H��t$�M����U�|
P t�E����M�TPR���E����M�|L t$�U����E�|T t�M����U�D
TP��넋M���   �´   R���E��]������������������������������������������������������������������������������������̋�U��Q�E���    ��   �M���   8���   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P�,�����M���   R�H0�����E���    t4�M���   �: u&j�E���   Q��+�����U���   P��/����j�M���   R�+����j�E���   Q�+�����U���    to�E���   �9 uaj�U���   -�   P�f+����j�M���   ��   R�L+����j�E���   ��   Q�2+����j�U���   P�+�����M���   ��t8�U���   ���    u&�M���   R�3����j�E���   Q��*�����E�    �	�U����U��}���   �E����M�|H��t:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP�n*�����M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!h0�j h�   h��j��������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ��)���������j�UR�)������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�{-�����}� t�E�P�.�����}� t�M��9 u�}�@�t�U�R�:�����E��]������������������������������������������̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    �,"���E��E��Hp#��t	�U��zl uDj�������E�    �D�P�M���lQ�`.�����E��E������   �j�)'��������!���Pl�U�}� u
j ��,�����E�M�d�    Y_^[��]������������������������������������������������������������U��WV�u�M�}�����;�v;���  ���   r�=<� tWV����;�^_u������   u������r)��$�Я�Ǻ   ��r����$���$����$�d���� �D�#ъ��F�G�F���G������r���$�Я�I #ъ��F���G������r���$�Я�#ъ���������r���$�Я�I ǯ���������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�Я��������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�l������$���I �Ǻ   ��r��+��$�p��$�l������̰�F#шG��������r�����$�l��I �F#шG�F���G������r�����$�l���F#шG�F�G�F���G�������V�������$�l��I  �(�0�8�@�H�P�c��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�l���|��������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�����M��)����U���   �P�� �  �M�M��,���E��]����������������������������̋�U��j �EP�����]�����������̋�U��h  �EP������]�������̋�U��h  �EP�����]�������̋�U��j�EP�����]����������̋�U��j�EP�q����]����������̋�U��j�EP�Q����]����������̋�U��j�EP�1����]����������̋�U��j�EP�����]����������̋�U��j�EP������]����������̋�U��h�   �EP������]�������̋�U��h�   �EP�����]�������̋�U��j�EP�����]����������̋�U��j�EP�q����]����������̋�U��j�EP�Q����]����������̋�U��j�EP�1����]����������̋�U��h  �EP�����]�������̋�U��h  �EP������]�������̋�U��hW  �EP������]�������̋�U��hW  �EP�����]�������̋�U��h  �EP�����]�������̋�U��h  �EP�n����]�������̋�U��j �EP�Q����]����������̋�U��j �EP�1����]����������̋�U���E=�   ���]������������̋�U��Qh  �EP��������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP�M������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Qh  �EP��������u�M��_t	�E�    ��E�   �E���]��������������������̋�U��Q3��} ���E��}� uh �j j$h��j�������u̃}� u-�e'���    j j$h��h`�h ��p!�����   ��U�d��3���]���������������������������������������̋�U��Q3��} ���E��}� uhP�j j-h��j�d������u̃}� u-��&���    j j-h��h0�hP��� �����   ��U�h��3���]���������������������������������������̋�U��Q3��} ���E��}� uh��j j6h��j��������u̃}� u-�%&���    j j6h��h��h���0 �����   ��U�`��3���]���������������������������������������̋�U����} t�} w�} u�} t	�E�    ��E�   �E��E��}� uh��j j?h��j� ������u̃}� u0�a%���    j j?h��hh�h���l�����   �<  �} t�U� 3��} ���E��}� uh4�j jDh��j�������u̃}� u0��$���    j jDh��hh�h4��������   ��   �} t�}t	�E�    ��E�   �U�U�}� uh��j jEh��j�������u̃}� u-�s$���    j jEh��hh�h���~�����   �Q�M����R���������M��} u3��,�U�;Ev�"   ��M����R�EP�MQ�%������]��������������������������������������������������������������������������������������������������������������������������������̋�U��d�]����̋�U��h�]����̋�U��`�]����̋�U����]����̋�U��j�hH�h9�d�    P��SVW���1E�3�P�E�d�    �=\� uEj������E�    �=\� u��   �\����\��E������   �j������ËM�d�    Y_^[��]����������������������������������������������̋�U��j�hh�h9�d�    P��SVW���1E�3�P�E�d�    j�������E�    �H   �E������   �j�K����ËM�d�    Y_^[��]�����������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �E�    �E�    j�0�����E�    �����E�j h�   h��h|�h<��E�P������P�����j h�   h��h|�h���M�Q�����P�{����j h�   h��h|�hx��U�R�����P�P�����?	���E��T�    �$������$���hx��������Eă}� t�M�����.  �=X� tj�X�P�S�����X�    h���8�����   �T�   ���k�<�M������t���k�<EЉE��B���t$�=P� t�E�   �P�+��k�<�U���E�    �E�    �E�Pj j?�M܋Rj�h��j �E�P����t�}� u�M܋�B? ��E܋� �U�Rj j?�E܋HQj�h �j �U�R����t�}� u�E܋H�A? �	�U܋B�  �E�   ��   �=X� t#�X�Q�U�R�2������u�E�   �   �=X� tj�X�P������h  h@�j�M�Q�
������P������X��=X� u	�E�   �Bj h  h��h|�h���U�R�E�P�q
������P�X�Q������P������U�R�\�����E�P�������M�Q������E������   �j�����Ã}� ��  j h-  h��h|�h��j�U�Rj@�E܋Q�����P������Uă��UċE����-u�Ũ��ŰEă��EċM�Q�����i�  �EЋU����+t�M����0|�E����9�Uă��U��ԋE����:��   �Uă��UċE�P�&����k�<EЉEЋM����0|�E����9�Uă��U��ߋE����:u<�Uă��UċE�P������EЉEЋM����0|�E����9�Uă��U��߃}� t�E��؉EЋM���Uԃ}� t8j h`  h��h|�hH�j�E�Pj@�M܋QR�H����P�K�����	�E܋H� �U�R�	�����E�P������M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���G����M�]���������������̋�U���]���M�]���������������̋�U���d���M�]���������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    j�z�����E�    �EP�T   ���E��E������   �j������ËE�M�d�    Y_^[��]��������������������������������̋�U����E�    j h.  h��h�h���E�P�	����P������}� u3��  �M�Q;�u�E�H;$���  �=T� �G  �@���uO�N�P�L�Q�J�R�H�Pj �D�Q�F�R�B�P�M�QRjj�g  ��,�G�N�P�L�Q�J�R�H�P�F�Qj j �B�R�E�HQj j�  ��,�����uO���P���Q���R���Pj ���Q���R���P�M�QRjj ��  ��,�G���P���Q���R���P���Qj j ���R�E�HQj j �}  ��,�   �E�   �E�   �E�   �E�   �U�zk}�E�   �E�   �E�
   �E�   j j j jj j �E�P�M�Q�U�BPjj�  ��,j j j jj j �M�Q�U�R�E�HQjj ��  ��,��;(�}K�E�H;�|�U�B;(�~3���   �M�Q;�~�E�H;(�}
�   �   �F�U�B;(�|�M�Q;�~
�   �   �E�H;(�~�U�B;�}3��e�M�Qk�<�E�ʋU�Bi�  �i��  �M��M�Q;�u�E�; �|	�   ��3����M�;,�}	�   ��3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �}�M  �E%  �yH���@��u�E��d   ����u#�El  ���  ����t�U�����E���M�����U��E����E��M��Fi�m  M��E���������E����d   ��+��E+  ���  ����D1�   ���U�U�;U�E+E�M��k�M�ȉM���U+U�Ek�E�E��}ud�M��  �yI���A��u�E��d   ����u#�El  ���  ����t�U�����E���M�����U�E�;E�~	�M����M��b�U��  �yJ���B��u�E��d   ����u#�El  ���  ����t�U�����E���M�����U�E�E��M�M �M��}u4�U����E$k�<E(k�<E,i��  E0� ��M���   �U��(��E$k�<E(k�<E,i��  E0�,�j h�  h��h8�hx��M�Q������P�A�����U�i��  ,��,�y �,� \&�,��(����(��+�=,� \&|�,��� \&�,��(����(��M�$�_^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�EP�M����3Ƀ} ���M�}� uh �j j4h��j��������u̃}� u=�g���    j j4h��hh�h ��r�����E�����M������E��  3��} ���E��}� uhL�j j5h��j��������u̃}� u=�����    j j5h��hh�hL��������E�����M��P���E��   �M�������z u"�EP�MQ��������EԍM�����E��x�b�U��E̍M��x���P�M�Q�������E��U���U�E��MȍM��N���P�U�R��������E��E���E�}� t�M�;M�t��U�+U��UЍM�����EЋ�]����������������������������������������������������������������������������������������������������������̋�U����E��M��U��E���E��A|�}�Z	�M��� �M��U��E��M��U���U��A|�}�Z	�E��� �E��}� t�M�;M�t��E�+E���]������������������������������̋�U����=�� ��   3��} ���E��}� uh �j jbh��j�e�������u̃}� u0�����    j jbh��h�h ���	���������   3҃} �U��}� uhL�j jch��j���������u̃}� u-�`���    j jch��h�hL��k	���������&�MQ�UR�d�������j �EP�MQ�������]������������������������������������������������������������������������̋�U��� V�E�    �E�E�3Ƀ} ���M�}� uh��j j6hx�j��������u̃}� u0�u���    j j6hx�h\�h��������   �u  j$h�   �EP�Q�����3Ƀ} ���M��}� uh4�j j:hx�j��������u̃}� u0�����    j j:hx�h\�h4�������   ��  �E��M��P�U�}�� |	�}�@W��s����    �   ��  �}�| 	�}��&A�v����    �   �  j h�3��E�P�M�Q�H�����F�E�E��F�j h�3�RP�$����M�+ȋE�M��E�E���������E����d   ��+ȋE�+  ���  ���D�j h�Q RP������M�+ȋE�M��E�}� }|�}� su�M����3��U�� �M��U�E���E�M��  �yI���A��u�E왹d   ����u�E�l  ���  ����u�U��Q �E�� �U��E�M����M��@�U��  �yJ���B��u�E왹d   ����u�E�l  ���  ����u	�U����U��E�M�Hj h�Q �U�R�E�P������M�A�U�B�j h�Q RP������M�+ȋE�M��E�}� t	�E�����E����E�   �	�M���M�U�E��M��;Q}��E���E�M�U�Q�E�M�U��@+��M�A�Uj h�Q �BP�
Q�F�������   ���E�Pj h  �M�Q�U�R�!����M�A�U�B�j h  RP������M�+ȋE�M��E�j j<�M�Q�U�R������M�A�U�Bk�<��M�+ȋE�U�
�E��@     3�^��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���������E��}� u3�� �EP�M�Q�x�����E��}� t3���E���]�������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� ������������������������������������������������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ���������������������������������������������̋�U����E�    �E�E�3Ƀ} ���M�}� uh��j j6h�j��������u̃}� u0�f���    j j6h�h��h���q�����   �2  j$h�   �EP�B�����3Ƀ} ���M�}� uh4�j j9h�j��������u̃}� u0�����    j j9h�h��h4��� �����   �  �E��M�}�@W��}����    �   �  �E��������E��U�iҀ��E�+E�M���F   �U��}�3�|[�E����E��M��3��M�}�3�|=�U����U��E�-�3��E�}� ��|�M����M��U�� ���U��	�E����E��M�U��Q�E����Q ���U�B�E�HiɀQ �U�+щU�}� t	�E�����E����E�   �	�E����E��M��U��E��;H}��U����U��E�M��H�U�E��M��R+��E�P�M����Q ������   ���E�P�E���  ���U�B�E�Hi�  �U�+щU�E���<   ���U�B�E�Hk�<�U�+ыE��M��A     3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �O����E��}� u�4���    3��N�E��xD u(h�   h��jj$�������E�M��U�QD�}� t�E��HD�M�������    3���E���]����������������������������������̋�U���������E��}� u3�� �EP�M�Q�^������E��}� t3���E���]�������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ���������������������������������������̋�U����} uh`�j jdhX�j�>�������u̋M�M��U�R�@������E��E��H��   u$���� 	   �U��B�� �M��A����G  �-�U��B��@t"�S��� "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6������ 9E�t������@9E�u�M�Q�[�������u�U�R��������E��H��  ��   �U��E��
+Hy!h��j h�   hX�j��������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�������E��q�}��t!�}��t�M����U���������U���E���E��H�� t7jj j �U�R�<������E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P�t������E�M�;M�t�U��B�� �M��A�����E%�   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hȥh9�d�    P���SVW���1E�3�P�E�d�    j��������E�    �E�x ��   ����M��E�����U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�������/�M�M��U�z uh`�j jXh��j�8�������u�랋M�QR��������E�@    �E������   �j������ËM�d�    Y_^[��]������������������������������������������������������������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �E�x �L  h (  h��h"�j �M��	Qj �v������E�}� u3��   �U�R�8������E��E��M����M���v�U�U���� u�M�M�� ��j�������E�    �U�z ��   j��������E܃}� ��   �E���P��������E؋M�U؉Q�}� t[j h�   h��hP�h���E�P�M���Q�U�BP�������P�>������M܋U�B��M܋U�B�A�M�U܉Q��E�P��������M�Q�M������E������   �j�������ËU�B�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    j�z������E�    �E�x ��   ����M��E�����U��U�}� tY�E�M�;Qu�E��M�Q�P�E�P�������2�M�M��U�z u!h`�j h�   h��j���������u�뛋M�QR��������E�@    �E������   �j�C�����ËM�d�    Y_^[��]���������������������������������������������������������������������̋�U���E��u	� (  f�M�URh��h"��EP�MQ�UR�>�����]���������������������̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    �E�x �a  j��������E�    �M�y �*  h (  j �U��	Rj �W������E�}� u"�E�    j��E�Ph���������E��  �M�Q�Y������E��U��E����E���v�M�M���� u�E�E��  ��j��������E܃}� ��   �E�    �M���Q�������E؃}� taj h4  h��h�h���U�R�E���P�M�Q�A�����P�������U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P�������M�Q�������E������   �j�������ËU�B�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������̋�U��j�hH�h9�d�    P���SVW���1E�3�P�E�d�    j�������E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P�g������M�Q�[��������E������   �j�������ËM�d�    Y_^[��]�����������������������������������������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�������������������������������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    �E�    j�������E�    �E�   �	�E����E��M�; 	��   �U����<� t|�M�������H��   t"�U�����Q����������t	�U���U�}�|=�E�������� R��j�E������R�������E������    �Y����E������   �j�������ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������̋�U����E�    �E�    �	�E����E��}�$}Z�M��<�D�uK�U�k����E���@��M����M�h�  �U���@�P����u�M���@�    3��뗸   ��]��������������������������������������̋�U����E�    �	�E����E��}�$}O�M��<�@� t@�U��<�D�t3�E���@��M��U�R��j�E�P��������M���@�    ��E�    �	�U����U��}�$}3�E��<�@� t$�M��<�D�u�U���@��E�M�Q��뾋�]��������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E�   �=l� u�+���j������h�   �������E�<�@� t
�   �   h  hP�jj�v������E�}� u������    3��   j
�������E�    �M�<�@� uDh�  �U�R����u"j�E�P�g����������    �E�    ��M�U��@��j�E�P�6������E������   �j
������ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������̋�U��E�<�@� u�MQ�<�������u
j��������U��@�P��]�����������������̋�U��E��@�Q��]��������̋�U��EPj �<h�   ������]����������������̋�U��   ]����̋�U���0�    ]���������������̋�U���]��������̋�U����} |�}}	�E�   ��E�    �E��E��}� u"h8�j jqh��j�L�������u�d����}� u.�����    j jqh��h��h8�����������   �}�t�U���t	�E�    ��E�   �E�E�}� u"h��j jvh��j���������u������}� u+�)����    j jvh��h��h���4���������/�}�u�U������E�����M��U�E�����E���]������������������������������������������������������������������������������������������̋�U����} |�}}	�E�   ��E�    �E�E��}� u%h8�j h�   h��j��������u������}� u0�����    j h�   h��h��h8�������������c�}�u�U�����Q�E�����M��}�uj����U�����'�}�uj����M������U�E�����E���]��������������������������������������������������������������̋�U��Q���E��M���E���]������������������̋�U���]����̋�U��j�h��h9�d�    P���PP  �h������1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P������ƅ���� h�  j ������Q������3�f������h�  j ������P�t�����ƅЯ�� h�  j ��ѯ��Q�W������} |�}|����*  �E�    �}��   h��������   j h  h��h��h��j
h   ��п��R�EP�F�����P�,�����hX��D�} t�M�������
ǅ����D�������R�Dh8��D��п��P�Dh��D�!���ǅ���������=  �} ��   ǅ̯��    �I������ȯ���<����     �UR�EPh�  h   ��Я��Q�p�������̯����̯�� }*j h*  h��h��hةj"j������R�2����� �������ȯ�����̯�� }8j h-  h��h��h��hL�h   ��Я��R������P��������}uV�} tǅ����4��
ǅ�����j h2  h��h��hP�������Ph   ��п��Q�Q�����P������j h4  h��h��h����Я��Rh   ��п��P�K�����P�X������}u�M������t8j h9  h��h��h��h��h   ��п��P�������P������j h:  h��h��h(�h�h   ��п��Q�������P��������} ��   ǅį��    �Z�����������M����     ��п��P�MQ�URh�h�  h   ������P�(�������į����į�� }*j hA  h��h��hةj"j������Q�7����� ��������������į�� }8j hD  h��h��h`�hL�h   ������P������P��������:j hH  h��h��h����п��Qh   ������R�v�����P������ǅ����    ǅ����    j�������Ph   ������Q������R�������������j hM  h��h��hH�j"j������P�F����� ������ t8j hO  h��h��h`�h��h   ������Q������P�������=,� u�=(� �#  ǅ����    ǅ����    j�+������E�   �,���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un�(���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j������Ã����� �D  �=� t?ǅ����    ������R������P�MQ������tǅ����   ������������������ ��   �E������t>�U�<����t1j ������P������Q������P������R�E����Q�@�U������t������Q�D�U������twƅп�� �} t9j h�  h��h��h��j
h   ��п��Q�UR�������P��������Я��P�MQ�U��ҍ�п��#�R�MQ�UR�Z������������E������   ��}uh����Ë������M�d�    Y_^[�M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hئh9�d�    P���\�  �8������1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q�~�����3�f������h�  j ������P�_�����ƅ���� h�  j ������Q�B�����3�f��Џ��h�  j ��ҏ��P�#������} |�}|����.  �E�    �}��   h��������   j h�  h��h0h�j
h   ��Я��Q�UR�N�����P�������hp�L�} t�E������
ǅ���H�����Q�Lh4�L��Я��R�Lh0�L�����ǅ���������A  �} ��   ����� ��ȏ�������     �MQ�URh�  h   ��Џ��P���������̏����̏�� }*j h  h��h0hةj"j�����Q������ ������ȏ�����̏�� }8j h  h��h0hxh��h   ��Џ��P�8�����P��������}uV�} tǅ���D�
ǅ���j h  h��h0hH �����Qh   ��Я��R�������P�h�����j h  h��h0h����Џ��Ph   ��Я��Q������P�.������}u�U������t8j h  h��h0h��hx�h   ��Я��Q�������P�������j h  h��h0h �h0h   ��Я��R������P�������} ��   ǅď��    �0���� �������#����     ��Я��Q�UR�EPh�h   h   ������Q��������ď����ď�� }*j h  h��h0hةj"j������R������ �������������ď�� }8j h  h��h0h �h��h   ������R�=�����P��������:j h"  h��h0h����Я��Ph   ������Q������P������ǅ����    j h(  h��h0h��j"jj�������Rh   ������Pj �������P�7����� ������������ t8j h*  h��h0h �h��h   ������Q������P��������=,� u�=(� �#  ǅ����    ǅ����    j�������E�   �,���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un�(���������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j������Ã����� �g  �=� t?ǅ����    ������R������P�MQ������t������������ǅ����   ������ �  �E�������[  �U�<�����J  �E����Q������������t�Jj ������R������P�������P������Q�U����P�H��t��   ����t��   ǅ���    j h{  h��h0h�j"jj�������Qh   �����R�����P�#�����P�t����� ���������� t>�����Pt5j ������Q������R�$�������P������P�M����R�@�@����� v������������j ������Q�����R�����P�M����R�@�E������t������R�L�E������ty3�f��Я���} t9j h�  h��h0h�j
h   ��Я��P�MQ�������P�~�������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ詾�����������E������   ��}uh����Ë������M�d�    Y_^[�M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�@��M�D��U�H��E�L�]�����������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �}t�}u�T  �}t�}t�}t�}t
�}�F  j �I������E�    �}t�}u=�=P� u4jh`�P��u�P�   ������	����0�E�   �E�E̋M̃��M̃}���   �U���@
�$�,
�@�Q�l�E�}t�UR���@��r�D�P�l�E�}t�MQ���D��L�H�R�l�E�}t�EP���H��%�L�Q�l�E�}t�UR���L��E������   �j ������Ã}� t��   ��   �}t�}t�}t��   �N����E؃}� u��   �E؁x\��uLhY  h(j�8�Q臸�����EȋU؋EȉB\�}� t�8�Qh���U؋B\P���������j�M؋Q\R�EP�5  ���E��}� u�L�M��Q�U�}t5�E��H;Mu*�U��E�B�M����M��<�k��E�P\9U�r��ˋE��   �M�MċUă��Uă}�w�E���`
�$�X
����x3�t	�E�   ��E�    �E��EЃ}� u!h�j h�  hhj虽������u̃}� u.������    j h�  hhhXh���������������M�d�    Y_^[��]Ë��;�` �I �	�	     ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    j ��������E�    �} u�E�@��E܋Q�l�E��E�   ��E�D��U܋P�l�E��E�   �}� t�}�t
�/����M܉�E������   �j ������Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������̋�U��j�hH�h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U���t�$�\�E�@��MЋ�U�E؃��E��  �E�D��MЋ�U�E؃��E���   �E�H��MЋ�U�E؃��E���   �E�L��MЋ�U�E؃��E��   萵���E��}� u�����  �M��Q\R�EP��  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!h�j h�  hhj蝹������u̃}� u1������    j h�  hhhdh�����������4  �E�P�l�E�}�u3��  �}� uj軻���}� t
j �K������E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<�0��M��	�Uԃ��Uԡ0�4�9E�}�M�k��U��B\�D    ���
�N����MЉ�E������   ��}� t
j �!�����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]Ë��^$A� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M��Q;Ut�E����E��<�k�M9M�s�ً<�k�U9U�s�E��H;Mu�E���3���]������������������������������������̋�U��H�P�l]�������������̋�U���ɾ����d]�����������������̋�U��詾����`]�����������������̋�U���@���3ŉE��E�    �׻���E��E�    �E�    �E�    �=X� ��   h�� �Eԃ}� u3��  h��E�P�T�E��}� u3��  �M�Q���X�h��U�R�TP���\�h��E�P�TP���`�h��M�Q�T�E��U�R���h��=h� tht�E�P�TP���d��d�;M�th�h�;U�t]�d�P�l�EЋh�Q�l�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�\�;M�t�\�R�l�Eȃ}� t�UȉE�}� t*�`�;E�t �`�Q�l�Eă}� t
�U�R�UĉE�X�P�l�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��Ю����]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� u!ht�j h�   hHj�;�������u̃}� u1�����    j h�   hHh0ht�����������Z  3Ƀ} ���M̃}� u!hj h�   hHj�Ѳ������u̃}� u1�2����    j h�   hHh0h�:����������   �E�E��M��AB   �U�E�B�M�U��E��@����M�Qj �UR�E�P�������E��} u�E��   �M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj ��������EċE�H���M��U�E��B�}� |!�M�� 3�%�   �E��M����E���M�Qj �������E��E���]��������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ��������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ蜸������]����������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR茻������]������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ��������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�ڷ������]��������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�ʺ������]����������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�?�������]��������������������̋�U��Q�E�E��M�Q�UR��������]����������������̋�U��Q�E�E��M�Q�UR��������]����������������̋�U��Q�E�E��M�Q�UR�EP�װ������]������������̋�U��Q�E�E��M�Q�UR�EP�=�������]������������̋�U����} u3��k  3��} ���E��}� uh �j j7hj�U�������u̃}� u0�����    j j7hh�h ���������   �  �} t�U;U��   �EPj �MQ聮����3҃} �U��}� uhL�j j=hj�˭������u̃}� u-�,����    j j=hh�hL��7������   �~�M;M҃��U�uh�j j>hj�j�������u̃}� u-������ "   j j>hh�h��־�����"   ��   ��MQ�UR�EP�v�����3���]������������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M���E����E���t��E�+E������]����������������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�j jh��j��������u̃}� u0�}����    j jh��h�h�舽�����   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E�M���Qh�   �U��R�	�����3��} ���E��}� uhL�j jh��j�S�������u̃}� u0�����    j jh��h�hL�迼�����   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P� ���������t3�t	�E�   ��E�    �E܉E�}� uh��j jh��j�3�������u̃}� u-����� "   j jh��h�h��蟻�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9��s����U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR������3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ����������������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]���������������������������������̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�������������������������������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    �e��E�   �E�    �E�P�E�������u�E�    �E������E��   �M+M�M܋U�R�E�P�Q������E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]������������������������������������������������������������������������������̋�U��E�p�]�����������������̋�U��Qj��������p�P�l�E��MQ���p�j�S������E���]�����������������̋�U��} th�j jWhj�q�������u�j �>�����]���������������������������̋�U��p�P�l]�������������̋�U��Q�p�P�l�E��}� t�MQ�U�����u3���   ��]��������������������������̋�U��Q�E�    �}�wC�EP�������E��}� t�*�=�� u�����    ��MQ�v�������u����UR�`������߻���    3���}� u�ʻ���    �E���]���������������������������������������̋�U��Q�=l� u�n���j������h�   �Ħ�����} t�E�E���E�   �M�Qj �l�R�T��]�������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �} t�}t	�E�    ��E�   �EԉE܃}� uhЧj jahX�j�B�������u̃}� u.裺���    j jahX�h�hЧ讴��������h  3҃} �U؃}� uh��j jbhX�j�ޢ������u̃}� u.�?����    j jbhX�h�h���J���������  j輣�����E�    �,��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���MЋU�EЉB�MЉM��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�,�j�U�R�)������43�uh��j jhX�j�ӡ������u��E������3����    ��   �}� tu�U�B���E̋M�ỦQ�ẺE��M�;,�tM�U�z t�E�H�U���M��E�H�J�U��    �E�,��H�,��E��M�,��h�   hL�jj�������E�}� u�E�����肸���    �L�U��    �E�,��H�=,� t�,��E��M��A   �E�   �U�E�B�M�,��E������   �j�K�����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP肟�����E��E�    �E���]�����������������̋�U��EP�MQ�UR�EP�MQ�UR肭����]���������̋�U��P  �.������3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �P��u8j h<  hX�h�	h�	hd	h  ������Q�G�����P舩�����������U��E�P財������@v]�M�Q衡�����U��D��E�j hE  hX�h�	hH�j���Q�U�������+й  +�Q�U�R�A�����P�������} t'�EP�>�������@v�MQ�-������U�DÉE�������������r����     �}uǅ������
ǅ����k��U���t�M�������
ǅ����k��U���t�}uǅ������
ǅ����k��M���tǅ������
ǅ����k��} t�E�������
ǅ����k��} tǅ������
ǅ����k��} t�M�������
ǅ����k��} tǅ������
ǅ����k��}� t�U��������'�} t�E�������
ǅ����k��������������}� tǅ������
ǅ����k��} tǅ������
ǅ����k�������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U���Ph8h�  h   ������Q衞����D�E�}� }*j h`  hX�h�	hةj"j�k����R趗���� �[�����������}� }8j he  hX�h�	h`�hL�h   ������R�4�����P�u�����h  h������P������������������uj�	�����j����������u�   �3��M�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���V3��} ���E�}� uh�
j jHhP
j��������u̃}� u-�r����    j jHhP
h,
h�
�}�����3��   �}�v�?����    3��~�} u�E   �URj �l�P�\�E��MQ�URj�l�P�X�E��}� u:�}� @  w�M;M�w�x   ��t�U�U����P�{�������輰���0�E�^��]����������������������������������������������������������������������������̋�U����E�����j j�E�Pj �l�Q�`��t�}�u	�E�   ��E�    �E���]�������������������������̋�U���V�E�E��} u�MQ�$�������   �} u�UR�w�����3��   �E�    �}�w)�} u�E   �EP�MQj �l�R�X�E���EP������耯���    3��e�}� u	�=�� u%�}� t���P���������I����0�E��1�MQ貤������u��P�۟�����������03���J���^��]����������������������������������������������������������������������̋�U��QV�E�    �} u�4�EPj �l�Q�d�E��}� u��P�=��������~����0^��]���������������������������������̋�U��Q�E�����j j �l�P����u�E������E���]�����������������̋�U���̘��]����̋�U���<�E�    3��E؉E܉E��E�E�E�E��MԉM�3҃} �UЃ}� uht�j jih j�>�������u̃}� u.蟭���    j jih h�
ht�誧��������  3Ƀ} ���M̃}� uhj jnh j�ڕ������u̃}� u.�;����    j jnh h�
h�F���������   �E�E��M��A����U��BB   �E�M�H�U�E��M�Qj �UR�E�P�������E��} u�E��Q�M�Q���UȋE�MȉH�}� |"�U��  3Ɂ��   �MċU����M���U�Rj ��������EċE���]��������������������������������������������������������������������������������������������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�a�������]������������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ蒨������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�P�������]��������������������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR��������]������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�=�������]����������������̋�U��Q�E�E��M�Qj �UR�EP�MQ衧������]����������������������̋�U��Q�E�E��M�Q�UR�EP�MQ�UR�_�������]��������������������̋�U��Q�E�E��M�Q�UR��������]����������������̋�U��Q�E�E��M�Q�UR胍������]����������������̋�U��Q�E�E��M�Q�UR�EP�;�������]������������̋�U��Q�E�E��M�Q�UR�EP耟������]������������̋�U��E��=   vh�j j8hxj��������u̋UR�EPj 見����]����������������������������̋�U����EP�M������M����   vh�j jDhxj�z�������u̃}�|5�}�   ,�M��ΐ��� ���   �U�Q#E�E�M��>����E��1�'�M�袐������   �B�#E�E�M������E���M�������]��������������������������������������������������̋�U���(�EP�M�蟚���}�|6�}�   -�M���������   �E�B#M�M��M�芨���E��   �M�����P�U�����   R赑������t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M�藏��� �HQ�M�艏����BP�M�Q�U�R�E�Pj�M��m���P�_����� ��u�E�    �M��ާ���E���M�#M�M؍M��ǧ���E؋�]������������������������������������������������������������������������������̋�U��=�� u�E���A#E��j �UR�EP�F�����]��������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E������E�    j���������u����C  j�������E�    �E�    �	�E���E�}�@��  �M�<��� �#  �U�����E��	�M؃�@�M؋U����   9E���   �M��Q����   �E؃x uaj
�_������E�   �M؃y u.h�  �U؃�R����u	�E�   ��E؋H���U؉J�E�    �   �j
莛����Ã}� u+�E؃�P���M��Q��t�E؃�P���4����}� u-�M��A�U�������E����M�U�+�����E��������}��t��   ��   h�   h,jj@j ��������E؃}� ��   �E�M؉����h��� �h��	�E؃�@�E؋M������   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃��������D�U�R��������u�E������������E������   �j�6�����ËE܋M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} ��   �E;h���   �M���U���������<�um�=��uB�M�M��}� t�}�t�}�t�(�URj��h��EPj��h��MQj��h�U���E���������U�3���艢��� 	   �5����     �����]�����������������������������������������������������������̋�U��Q�} ��   �E;h���   �M���U���������L����   �U���E���������<�th�=��u<�U�U��}� t�}�t�}�t�"j j��h�j j��h�
j j��h�E���M�������������3����j���� 	   �����     �����]������������������������������������������������������������̋�U����}�u躏���     ������ 	   ����2  �} |�E;h�s	�E�   ��E�    �M�M��}� u!h8�j h;  h�j�0�������u̃}� u<�H����     膠��� 	   j h;  h�hhh8�莚��������   �E���M���������D
������؉E�u!h��j h<  h�j褈������u̃}� u9輎���     ������ 	   j h<  h�hhh�������������U���E�����������]����������������������������������������������������������������������������������������������̋�U��j�hاh9�d�    P���SVW���1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP���E��}� u��P�l���������q  �}�u�M��@�M���}�u
�U���U��)����E؃}��u�|����    �(����     ����#  �E�    �EP�M�Q��������U���U�E����M؃��������E�D
�M����U؃��������L$�ဋU����E؃��������L$�E����M؃��������D
$$�M����U؃��������D$�E�   �E������   �K�}� u8�U����E؃��������T����E����M؃��������T�M�Q�J�����Ã}� t�U؉U���E������EԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E���M��������M��E�   �U��z u_j
�������E�    �E��x u,h�  �M���Q����u�E�    �U��B���M��A�E������   �j
������Ã}� t!�U���E���������TR���E�M�d�    Y_^[��]��������������������������������������������������������������������������̋�U��E���M���������D
P��]������������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �}�u�ٚ��� 	   ����  �} |�E;h�s	�E�   ��E�    �M؉M��}� uh�j j,h`j��������u̃}� u.�u���� 	   j j,h`hHh�耔��������;  �E���M���������D
������؉E�uhj j-h`j虂������u̃}� u.������ 	   j j-h`hHh�����������   �UR�~�����E�    �E���M���������D
��t;�MQ� �����P�l��u���E���E�    �}� u�>�����U��^���� 	   �E�����3�uh��j jEh`j�Á������u��E������   ��UR�~����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h8�h9�d�    P���SVW���1E�3�P�E�d�    �}�u������     �.���� 	   ����  �} |�E;h�s	�E�   ��E�    �M؉M��}� uh8�j jChpj�i�������u̃}� u9聆���     迗��� 	   j jChph`h8��ʑ��������/  �E���M���������D
������؉E�uh��j jDhpj��������u̃}� u9������     �9���� 	   j jDhph`h���D���������   �UR��{�����E�    �E���M���������D
��t�MQ�UR�EP�{�����E��?迖��� 	   �k����     �E�����3�uh��j jOhpj�������u��E������   ��EP�\{����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U�츐<  �>}�����3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uhpj jmhpj��}������u̃}� u9�����     �?����    j jmhphLhp�J���������
  �E���M���������D
$�����E��M���t	�U���uo�E��������E�uh$j juhpj�G}������u̃}� u9�_����     蝔���    j juhphLh$討���������	  �U���E���������T�� tjj j �EP�}�����MQ��������td�U���E���������T��   tA�����EԋEԋHl3҃y �U�E�P�M���U���������Q�t�E�}� ��  �}� t�U�����  �p�E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M���������|
8 ��   �E���M���������D
4P�v������u!h�j h�   hpj�{������u̋U���E���������T4�U��EЊ�M��U���E���������D8    j�U�R�E�P�z�������u�  �   �M��R�u��������   �E�+E�M+ȃ�v'j�U�R�E�P�Pz�������u�O  �MЃ��M��K�U���E���������UЊ�T4�E���M���������D
8   �E����E���  �j�M�Q�U�R��y�������u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R���Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M���������
P�@��t�M�+MM�M��U�;U�}�  ����E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M���������
P�@��t!�M�;M�}�   �U���U�E����E�����E��   �   �M���t	�U���u{�E�P�/��������U�;�u�E����E�����E��R�}� tG�E�   �   f�M��U�R���������M�;�u�U����U��E���E�����E���t�����  �M���U���������L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E���������R�@��t �E�E��E�������������+�9M�}�����E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U���������Q�@��t �U�U��U�������������+�9E�}�����E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  ����t�����t��� u���E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E���������R�@��t��p���E���p�������E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U���������Q�@��t�E�    �U��U��	���E�}� ��   �}� t0�}�u����� 	   �y���M���U�R�q��������V�L�E���M���������D
��@t�M���u3��%�貊���    �^y���     ������E�+E�M�3���m����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hX�h9�d�    P���SVW���1E�3�P�E�d�    �}�u�0v���     �n���� 	   ����(  �} |�E;h�s	�E�   ��E�    �MԉM��}� uh8�j jTh�j�o������u̃}� u9��u���     ������ 	   j jTh�h�h8��
���������  �E���M���������D
������؉E�uh��j jUh�j�#o������u̃}� u9�;u���     �y���� 	   j jUh�h�h��脀��������  ����;U����E�uh�j jVh�j�n������u̃}� u9��t���     �
����    j jVh�h�h�����������   �UR�j�����E�    �E���M���������D
��t�MQ�UR�EP�si�����E��?萅��� 	   �<t���     �E�����3�uh��j jah�j��m������u��E������   ��EP�-j����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���tV�E������E�E��}�u�s���     �J���� 	   ����	  �} |�M;h�s	�E�   ��E�    �U��U��}� u!h8�j h�   h�j�l������u̃}� u<�r���     �؃��� 	   j h�   h�h�h8���}��������y  �M���U���������L������ىM�u!h��j h�   h�j��k������u̃}� u<�r���     �L���� 	   j h�   h�h�h���T}���������  ����;EɃ��M�u!h�j h�   h�j�k������u̃}� u<�q���     �ׂ���    j h�   h�h�h���|��������x  �E�    �} t �E���M���������D
��t3��D  3Ƀ} ���M��}� u!hxj h�   h�j��j������u̃}� u<��p���     �.����    j h�   h�h�hx�6|���������  �E���M���������D
$�����E�M�M��}�t�}��  �  �U����҃��U�u!h$j h�   h�j�'j������u̃}� u<�?p���     �}����    j h�   h�h�h$�{��������  �M���s	�E�   ��U��U��E��Eh�   h@j�MQ�c�����Eԃ}� u�
����    �o���    ����  jj j �UR�0j�����M���u���������D1(�T1,�   �U����҃��U�u!h$j h�   h�j�i������u̃}� u<�5o���     �s����    j h�   h�h�h$�{z��������  �M����M�U�UԋEԉEȋM���U���������L��H��  �U���E���������T��
�r  �} �h  �E���M���������EȊL
��Uȃ��UȋẼ��E̋M���M�U���E���������D
�U���  �E���M���������D
%��
��   �} ��   �M���U���������MȊT%��Eȃ��EȋM̃��M̋U���U�E���M���������D
%
�E��u{�M���U���������L&��
t[�} tU�U���E���������UȊD&��Mȃ��MȋŨ��ŰE���E�M���U���������D&
j �M�Q�UR�E�P�M���U���������Q�x��t�}� |�U�;Uv^���E܃}�u#�$~��� 	   ��l���M܉�E������  �,�}�mu�E�    �  ��U�R�d�����E������|  �E�E�E̋M���U���������L��   �L  �U����  �}� tE�E����
u:�U���E���������T���E���M���������T�8�M���U���������L����U���E���������L�EԉE؋M؉M��U�U�9U��9  �E������   �U���E���������T��@u:�E���M���������D
���M���U���������D��U؋E���
�U؃��U؋E����E��  �  �M����t!�E؋M����E؃��E؋M����M��y  �ŰEԍL�9M�sG�U��B��
u�M����M��U��
�E؃��E���M؋U����M؃��M؋U����U��#  �E����E��E�    j �M�Qj�U�R�E���M���������
P�x��u	���E܃}� u�}� u�M���U؃��U��   �E���M���������D
��HtH�M��
u�U��
�E؃��E��,�M���U؃��U؋E���M���������E�D
�R�M�;M�u�U��
u�E�� 
�M؃��M��0jj�j��UR�:d�����E��U��E��
t�M���U؃��U������E�+EԉE��M����  �}� ��  �U؃��U؋E����   u�U؃��U��O  �E�   �E��������u"�}��E�;E�r�M؃��M؋U����U��͋E�������U��}� u�,z��� *   �E������  �E���;E�u�M�M��M���   �U���E���������T��H��   �E���M���������E؊ �D
�M؃��M؃}�|(�U���E���������U؊�T%�E؃��E؃}�u(�M���U���������M؊	�L&�U؃��U؋E�+E��E��j�E��ؙRP�MQ�b�����E��UċU�+UԉŰE���P�MQ�U�R�E�Pj h��  ��Ẽ}� u��P�_�����E������  �M�+M�3�9M��E���M���������T0�M���M��S  �}� tE�U����
u:�M���U���������L���U���E���������L�8�E���M���������D
����M���U���������D�UԉU��E��EЋM�M�9M���  �U������   �M���U���������L��@u:�U���E���������T���E���M���������T��M��U�f�f��M����M��UЃ��U��   �  �E����t#�U��E�f�f�
�U����U��EЃ��E���  �M̋UԍD
�9E�sN�M��Q��
u�EЃ��Eй
   �U�f�
�E����E���M��U�f�f��M����M��UЃ��U��  �EЃ��E��E�    j �M�Qj�U�R�E���M���������
P�x��u	���E܃}� u�}� u�   �U�f�
�E����E��  �M���U���������L��H��   �U��
u�
   �M�f��U����U��|�E�E��   �U�f�
�E����E��M���U���������M��	�L�U����U��E���M���������E�� �D
%�M���U���������D&
�\�M�;M�u�U��
u�
   �M�f��U����U��5jj�j��EP��^�����E��U��M��
t�   �E�f��M����M��E����U�+UԉŰE�;Et�M�Q�{t�����}��u�ỦU���E�E��E�^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} uh`�j j.hj�Y������u̋��������U�U�j:h�jh   �zS�����E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]��������������������������������������������������������������̋�U��j�hx�h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E������E�    3��} ���EЃ}� uh j jhh�j�sX������u̃}� u.��o���    j jhh�h�h ��i���������   �U�UԋEԃ��EԋMԋQ��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q��  ���E��E������   �Q�}� tJ�}� t8�U����E؃��������T����E����M؃��������T�M�Q��S����Ã}� t��n���U�������E؋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E�    3��} ���E܃}� u!h�j h�   h�j�V������u̃}� u3��m���    j h�   h�h�h��h�����   �  �U�����3��} ���E؃}� u!h j h�   h�j�)V������u̃}� u3�m���    j h�   h�h�h �g�����   �  �} to�U�������҃��U�u!h(j h�   h�j�U������u̃}� u3�m���    j h�   h�h�h(�g�����   �   �E�    �MQ�UR�EP�MQ�UR�EP�M�Q�)  ���E��E������   �[�}� tT�}� t@�U����M����������L����U����U����������L�M�R�BQ����Ã}� t	�E� �����E�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �E�    �E� �E�    �E�   �E�    �E%�   t�E�    �E���E�   �E� j h�   h�h�h��M�Q�$b����P�~^�����U�� �  u/�E% @ t�M��ɀ   �M���}� �  t�U��ʀ   �U��E���E�t�}�t�}�t6�@�E�   ���   �M��t�U��   t	�E�   ���E�   @�   �E�   ��   �=Y���     �E� ����3�t	�E�   ��E�    �U��U��}� u!h�j h	  h�j��R������u̃}� u3�+j���    j h	  h�h�h��3d�����   �  �M�M��U����U��}�pw_�E������$����E�    ��   �E�   ��   �E�   �   �E�   �   �}�   �u	�E�   ��E�    �   �;X���     �U�����3�t	�E�   ��E�    �M��M��}� u!h<j h,  h�j��Q������u̃}� u3�)i���    j h,  h�h�h<�1c�����   �  �E%   �E��}�   7�}�   tK�}�   �}�   t]�}� t3�}�   t6�d�}�   tO�Y�}�   t,�}�   t/�}�   t�<�E�   �   �E�   �   �E�   �   �E�   �   �E�   �   �	W���     �M�����3�t	�E�   ��E�    �E��E��}� u!h�j hN  h�j�P������u̃}� u3��g���    j hN  h�h�h���a�����   �  �E�   �U��   t�����#E%�   u�E�   �M��@t �U��   �U�E�   �E��M���M�U��   t�E�   �E�M�� t�U��   �U���E��t�M��   �M���h���U��E�8�u+��U���     �M������g���    �g��� �
  �U�   j �E�P�M�Q�U�R�E�P�M�Q�UR�|�E��}���  �E�%   �=   ���   �M����   �U�������U�j �E�P�M�Q�U�R�E�P�M�Q�UR�|�E��}��u^�E����U����������T����E����E� ���������T��P��L�����f����U���	  �^�E����U����������T����E����E� ���������T��P�tL�����e����U��g	  �E�P���E�}� ��   �E�    �M����E����������D
����M����M�	���������D
���E��E�P��K�����M�Q���}� u�*e���    �e����U���  �}�u�E���@�E���}�u
�M����M��U�R�E�Q�H�����U����U��E����U����������U��T�E����U����������T$�​E����E� ���������T$�U���H��   �E�%�   ��   �M����   jj��U�P�P�����Eă}��u/��R���8�   t�M�R�6T�����d��� �E��  �   �E� j�M�Q�U�P��G������u?�Mσ�u6�EęRP�U�P�'W�������u�M�R��S�����c��� �E��_  j j �M�R�	P�����Eă}��u�E�Q�S�����|c����U��'  �E�%�   �;  �M�� @ u'�Uȁ� @ u�E @  �E��Mȁ� @ M�M�U�� @ u!h�j h&  h�j�K������u̋M�� @ ��|�����|���   2��|���   ti��|��� @  t@��|���   t:��|��� @ t.�M��|��� @ t7��|���   t1��|��� @ t%�'�E� �!�U��  ��  u�E��
�E���E��E%   �5  �E�    �E�    �E�    �M���@��  �U���   ���x�����x���   @t-��x���   �t��x���   ���   �  �E�   �  �EЉ�t�����t�������t�����t�����   ��t����$�0�jj j �E�Q��J������l�����p�����l����p���tPj j j �E�Q��J������d�����h�����d���#�h������u�E�Q�qQ�����Oa����U���  ��E�   ��   �EЉ�`�����`�������`�����`�����   ��`����$�D�jj j �E�Q�BJ������X�����\�����X����\���tWj j j �E�Q�J������P�����T�����P���#�T������u�E�Q�P�����`����U��>  �E�   ��E�   ��E�   �}� ��  j�E�P�M�R�+D�����E��}� ~2�}�u,3�u!htj h�  h�j�H������u��E�    �U���L�����L����t��L���t=��L���t"��   �E�Q��O������_����U��  �}�﻿ u	�E���   �E�%��  =��  uJ�M�R�O����3�u!h�j h�  h�j�H������u��x_���    �E�   �  �U�����  ����  u>j j�E�Q�K�����Eă}��u�U�P�IO�����'_����M���  �E��8j j �U�P�vK�����Eă}��u�M�R�O������^��� �E��  �}� ��   �E�    �E�    �E�    �MH�����H���t��H���t��E���  �E�   ��E�﻿ �E�   �U�;U�~U�E�    �E�+E�P�M��T�R�E�Q�F�����E��}��u�U�P�_N�����=^����M���  �U�U��U�룋E����U����������U���D$$�
M����M�	���������D
$�E%   ����؋M����M�	��������$���L
$��
ȋU����U����������L$�M���HuH�U��t@�E����U����������T�� �E����E� ���������T�U���   ���   ���   �E����   �M�Q���U�������U��E�   j �E�P�M�Q�U�R�E�P�M�Q�UR�|�E��}��uk��P�zC�����E����U����������T����E����E� ���������T�U�P�>^�����t\����M��"� �U����M����������M���E���]Ë�uu'u3u?u]u �I �}�}%}%}�}o~o~�}�}o~�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR�I�����E�}� t	�E�������E��E�E��]������������������������������̋�U��j�EP�MQ�UR�EP�MQ�H����]�����������̋�U���HV�EP�M��I���} u�E�    �M��(W���E��d  �M��>���H�y u'�UR�EP�MQ�M�����E؍M���V���E��,  3҃} �U�}� uh�j j?h`j��>������u̃}� u=�!V���    j j?h`h<h��,P�����E�����M��}V���E��  3Ƀ} ���M��}� uh j j@h`j�M>������u̃}� u=�U���    j j@h`h<h �O�����E�����M��
V���E��F  �E�M���M���   �Uf�f�E��M���M�M��E=���P�E��L���	  �} u@3�f�U��M��=���@�M��D��t	�E�    �	�M��U�f�E�f�E��Y  �M���u3�f�E��   �M����U��f�M��M���M�u��M��<���P�B;�|2�u��M��<���H�Q;��M��<���@�H�U��f�U��G�u��M��d<���@�H;�|0�u��M��M<���P�B;��M��:<���H�Q�E��f�E��D�M��<���H�U��D��t�M��<���H�U���  �E���M��M�f�U�f�U��Ef�f�M��U���U�M���;���@�M��T����   �} u3�f�E��  �M���M�U���u3�f�M��   �U����E��f�U��U���U�u��M��[;���@�H;�|2�u��M��D;���P�B;��M��1;���H�Q�E��f�E��G�u��M��;���H�Q;�|0�u��M���:���@�H;��M���:���P�B�M��f�M��D�M���:���P�E��L��t�M��:���P�E���  �M���U��U�f�E�f�E��M��U�;�t#�E��M�3�;��T��U̍M���R���E��3�E���u�E�    �M���R���E��������E�    �M��R���E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR��N����]�������������������̋�U���D�} u3���  �EP�M��C���M��8���H�y u'�UR�EP�MQ�I�����E܍M��Q���E��  3҃} �U�}� uh�j j>hj��8������u̃}� u=�2P���    j j>hh�h��=J�����E�����M��P���E��  3Ƀ} ���M��}� uh j j?hj�^8������u̃}� u=�O���    j j?hh�h ��I�����E�����M��P���E��  �E�M���M���s  �Uf�f�E��M���M�M��V7���P�E��L��t|�} u@3�f�U��M��17���@�M��D��t	�E�    �	�M��U�f�E�f�E��   �M���u	�E�    ��E����M�E��E���Ef�M�f�M��Uf�f�E��M���M�M��6���P�E��L��tM�} u3�f�U��?�E���E�M���u	�E�    ��E����M�E��E���Ef�M�f�M��U��E�;�t#�M��U�3�;����D ��EЍM��N���E��3�M���u�E�    �M��N���E���y����E�    �M��}N���Eȋ�]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR��C����]��������������������U��SVWUj j h��u�@��]_^[��]ËL$�A   �   t2�D$�H�3���/��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�u�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� �������������������������������������������������������������������������������������������̋�U����}�u�SK��� 	   3��   �} |�E;h�s	�E�   ��E�    �M��M��}� uh8�j j(h�j�3������u̃}� u*��J��� 	   j j(h�h�h8���D����3���E���M���������D
��@��]���������������������������������������������������̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uh�j jJhpj�2������u̃}� u0�J���    j jJhphPh��D�����   �\  �UR�M��8<���M���1��� �x ��   �M���   ~C�} t�} v�URj �EP�2�����I��� *   �}I����M؍M���I���E���  �} tw3�;U��؉E�uh��j j]hpj��1������u̃}� u=�+I��� "   j j]hphPh���6C�����E�"   �M��I���E��x  �U�E��} t	�M�   �E�    �M��YI���E��J  �=  �E�    �U�Rj �EP�MQj�URj �M��0��� �HQ���E��}� t
�}� ��   �}� ��   ����z��   �} t�} v�URj �EP�_1����3�t	�E�   ��E�    �U��U܃}� uhj j{hpj�0������u̃}� u:��G��� "   j j{hphPh�B�����E�"   �M��XH���E��L��G��� *   �G����MȍM��6H���E��*�} t�U�E���E�    �M��H���E���M��H����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�6����]��������������̋�U��� �E������EP�M���8���M��b.��P�MQ�M��T.������   P�MQ�U�R�J6�����E�}� u�E��E���E������M��M�M��F���E��]�����������������������������������������̋�U����E�����j �EP�<C��P�MQ�U�R��5�����E��}� u�E��E���E������E��]����������������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� ������������������������������������������̋�U���<  ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���6���E�    �D���E�3Ƀ} �������������� u!h�j h  h��j��,������u̃����� uF�;D���    j h  h��hTh��C>����ǅ��������M��D��������#  �E�������������Q��@��   ������P�x5�����������������t-�������t$����������������������������
ǅ�������������H$�����х�uV�������t-�������t$����������������������������
ǅ�������������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!h`�j h  h��j�h+������u̃����� uF��B���    j h  h��hTh`���<����ǅ��������M��C��������  3Ƀ} �������������� u!ht�j h  h��j��*������u̃����� uF�>B���    j h  h��hTht��F<����ǅ��������M��B��������&  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���  ������ �	  �������� |%��������x�������� ���������
ǅ����    ������������������k�	�������� ����������������   3�tǅ����   �
ǅ����    ������������������ u!h j ha  h��j�t)������u̃����� uF��@���    j ha  h��hTh ��:����ǅ��������M��(A��������  ��������������������  �������$� ��E�    �M��[(��P������R�(*��������   ������P�MQ������R�u  ���E��������U���U����������؉�|���u!hh�j h�  h��j�r(������u̃�|��� uF��?���    j h�  h��hThh���9����ǅ��������M��&@��������  ������R�EP������Q��  ����  �E�    �UЉUԋEԉE�M�M��E�    �E������E�    �  �������������������� ������������wK��������X��$�@��E����E��,�M����M��!�U����U���E��   �E��	�M����M��'  ��������*u(�EP�x<�����E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�<�����Ẽ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  �����������$�l��E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��P
  ��������������������A������������7�  ����������$����U���0  u�E�   �E��M���  tUǅx���    �UR��4����f������������Ph   ������Q�U�R�f=������x�����x��� t�E�   �&�EP��9����f��t�����t����������E�   �������U��W  �EP��9������p�����p��� t��p����y u� ��U��E�P�l'�����E��P�M���   t&��p����B�E���p�����+����E��E�   ��E�    ��p����B�E���p�����U���  �E�%0  u�M���   �M��}��uǅ��������	�Ủ�������������h����MQ��8�����E��U���  te�}� u���E��E�   �M���d�����h�����h�������h�����t��d������t��d�������d����ɋ�d���+M����M��[�}� u	� ��U��E���l�����h�����h�������h�����t��l������t��l�������l����ɋ�l���+E��E��  �MQ�8������`����2/������   3�tǅ����   �
ǅ����    ��������\�����\��� u!h�j h�  h��j�|"������u̃�\��� uF��9���    j h�  h��hTh���3����ǅ ��������M��0:���� �����  ��  �U��� t��`���f������f����`�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Bh�  h��j�Ú�]  R�J�����E��}� t�E��E��Ḿ�]  �M���Ẹ   �U���U�E�H��P���P�����T����M�� ��P�E�P�M�Q������R�E�P�M�Q��P���R�H�P�l�Ѓ��M���   t$�}� u�M��: ��P�U�R�T�P�l�Ѓ���������gu*�U���   u�M�� ��P�E�P�P�Q�l�Ѓ��U����-u�M���   �M��U����U��E�P�b#�����E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�&������@�����D����   �U���   t�EP��%������@�����D����   �M��� tB�U���@t�EP�4��������@�����D�����MQ�|4���������@�����D����=�U���@t�EP�V4�������@�����D�����MQ�;4����3҉�@�����D����E���@t@��D��� 7|	��@��� s,��@����ً�D����� �ډ�8�����<����E�   �E����@�����8�����D�����<����E�% �  u&�M���   u��8�����<����� ��8�����<����}� }	�E�   ��M�����M��}�   ~�E�   ��8����<���u�E�    �E��E��M̋Ũ��U̅���8����<���t{�E��RP��<���Q��8���R�}5����0��L����E��RP��<���P��8���Q��3����8�����<�����L���9~��L����������L����E���L�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅4����M���u������R�EP��4���Qj �K	  ���U�R������P�MQ�U�R�E�P�|	  ���M���t$�U���u������P�MQ��4���Rj0� 	  ���}� ��   �}� ��   ǅ���    �E���0����M܉�,�����,�����,�������,�������   ��0���f�f������������Pj�� ���Q��(���R�w4�����������0�������0�������� u	��(��� uǅ���������*�M�Q������R�EP��(���Q�� ���R�{  ���V�����E�P������Q�UR�E�P�M�Q�U  �������� |$�U���t������P�MQ��4���Rj ��  ���}� tj�E�P�m)�����E�    ����������� t������tǅ����    �
ǅ����   ���������������� u!h�j h�  h��j��������u̃���� uC�/2���    j h�  h��hTh��7,����ǅ���������M��2����������������������M��i2���������M�3������]ÍI {�w����l�x������������ �I '�ۡ���� ���3�s�M�ݢ��I�+�����F���=�Y�4�   	
�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�%�����E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����'  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tE�U�;U�u.�E�H��  ����ًU��  �����;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���(  ���3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T������ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    ��%����|���3Ƀ} ����0�����0��� u!h�j h  h��j�(������u̃�0��� uI�%���    j h  h��h�!h������ǅ ���������T�����%���� �����7  �E��,�����,����Q��@��   ��,���P��������(�����(����t-��(����t$��(�������(������������\����
ǅ\�������\����H$�����х�uV��(����t-��(����t$��(�������(������������X����
ǅX�������X����B$�� ���ȅ�tǅT���    �
ǅT���   ��T�����$�����$��� u!h`�j h  h��j�������u̃�$��� uI�$���    j h  h��h�!h`������ǅ����������T����a$���������T6  3Ƀ} ���� ����� ��� u!ht�j h  h��j�%������u̃� ��� uI�#���    j h  h��h�!ht������ǅ����������T�����#����������5  ǅL���    �E������ǅ@���    ���@�������@�����@����q5  ��@���u������ u�Z5  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Uǅ��������ǅ��������ǅp�������ǅ���������E���G�����G����E���E����1  ��L��� ��1  ��G����� |%��G�����x��G����� ����P����
ǅP���    ��P�����H�����H���k�	��8����� ����8�����8�����  �E���%��  �������u\j
��t���R�EP�������~9��t������$u+��@��� uh@  j ������P�
����ǅ����   �
ǅ����    �������)  j
��t���Q�UR���������������t������E��@��� ��   ������ |#��t������$u������d}ǅL���   �
ǅL���    ��L������������� u!h(!j hQ  h��j�B	������u̃���� uI� ���    j hQ  h��h�!h(!�����ǅ����������T����� ����������2  ������;�x���~��������H������x�����H�����H�����x����   ��8�����   3�tǅD���   �
ǅD���    ��D������������� u!h j h]  h��j�Z������u̃���� uI����    j h]  h��h�!h ������ǅ����������T���� ����������1  ��8�����@�����@�����.  ��@����$�����@��� u	������t��@���u�������u�.  ǅ����    ��T������P��G���R����������   ��L���P�MQ��G���R�9A  ���E���G����U���U��G�������؉����u!hh�j h�  h��j�&������u̃���� uI����    j h�  h��h�!hh������ǅ����������T���������������0  ��L���R�EP��G���Q�@  ���-  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �P-  ��G�����<�����<����� ��<�����<���wi��<��������$������������������D���������������3���������������"�������   ����������������������,  ��G�����*��  ������ u�EP�������������^  j
��t���Q�UR����������������t������E��@��� ��  ������ |#��t������$u������d}ǅ8���   �
ǅ8���    ��8������������� u!hp j h�  h��j��������u̃���� uI�[���    j h�  h��h�!hp �c����ǅ����������T�������������.  ������;�x���~��������4������x�����4�����4�����x����������������� uE��������Ǆ����   ����������G������������������������������   ������P��G���Qj��������������P���������؉����u!h�j h�  h��j��������u̃���� uI�$���    j h�  h��h�!h��,����ǅ����������T����w���������j-  �\*  �+������������������������Q�}���������������� }���������������������؉������������k�
��G����DЉ�������)  ǅd���    ��)  ��G�����*��  ������ u�UR��������d����^  j
��t���P�MQ����������p�����t������U��@��� ��  ��p��� |#��t������$u������d}ǅ0���   �
ǅ0���    ��0������������� u!hj h�  h��j�������u̃���� uI�w���    j h�  h��h�!h�����ǅ����������T��������������+  ��p���;�x���~��p�����,������x�����,�����,�����x�����p����������� uE��p�����Ǆ����   ��p�������G�����������p������������������   ������R��G���Pj��p�����������R�!	��������؉� ���u!hhj h�  h��j�� ������u̃� ��� uI�@���    j h�  h��h�!hh�H����ǅ����������T�������������*  �x'  �+��p�����������������������P�������d�����d��� }
ǅd����������d���k�
��G����DЉ�d����'  ��G�����(�����(�����I��(�����(���.�B  ��(��������$����U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅ8���    �*����"�������� �������������   �������%  ��G�����$�����$�����A��$�����$���7��"  ��$�����L��$����������0  u������   ��������������  �_  ǅ����    ������ u�UR�����f��<�����  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!hj h�  h��j���������u̃����� uI�!���    j h�  h��h�!h�)����ǅ����������T����t���������g'  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�����u!h`j h�  h��j��������u̃����� uI����    j h�  h��h�!h`�����ǅ����������T����d���������W&  �   �,��������������������������P�����f��<�����<���Qh   ��P���R������P����������������� t
ǅl���   �*  ������ u�MQ�����f��������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hj h�  h��j�n�������u̃����� uI�����    j h�  h��h�!h������ǅ����������T�������������%  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q���������؉�����u!h�j h�  h��j�^�������u̃����� uI����    j h�  h��h�!h�������ǅ����������T�������������$  �j  �,��������������������������R�����f��������������P���ǅ����   ��P����������  ������ u�UR��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hj h�  h��j�4�������u̃����� uI����    j h�  h��h�!h�
����ǅ����������T���������������"  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�c ��������؉�����u!h j h�  h��j�$�������u̃����� uI����    j h�  h��h�!h �	����ǅ����������T���������������!  �0  �+��������������������������P������������������ t�������y u#� �������������P�{������������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������a  ������%0  u��������   ��������d����uǅ���������d������������������������� u�MQ��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hj h6  h��j�4�������u̃����� uI����    j h6  h��h�!h�����ǅ����������T���������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�c���������؉�����u!h j h:  h��j�$�������u̃����� uI����    j h:  h��h�!h �����ǅ����������T���������������  �0  �+��������������������������R��	����������������%  tx������ u��������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������i������ u� �����������������������������������������t���������t���������������ɋ�����+������������  ������ u�UR��������������  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hj h�  h��j�/�������u̃����� uI�
���    j h�  h��h�!h�����ǅ����������T�����
����������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R�^���������؉�����u!h j h�  h��j��������u̃����� uI�}	���    j h�  h��h�!h �����ǅ����������T�����	����������  �+  �+��������������������������P���������������������   3�tǅ���   �
ǅ���    ����������������� u!h�j h�  h��j�>�������u̃����� uI����    j h�  h��h�!h������ǅ����������T���������������  �J  �������� t������f��L���f����������L����ǅl���   �  ǅh���   ��G����� ��G�����������@��������������  ��@��� ��  ������ |������d}ǅ���   �
ǅ���    ����������������� u!hj h�  h��j��������u̃����� uI�j���    j h�  h��h�!h�r����ǅ����������T�������������  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�H���������؉�����u!hxj h�  h��j�	�������u̃����� uI�g���    j h�  h��h�!hx�o ����ǅ����������T�������������  �  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��G�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Zh�  h��j��d�����]  R�
����������������� t ��������������d�����]  ��P����
ǅd����   ������ u#�U���U�E�H��P��������������  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u!hj h  h��j�`�������u̃����� uI����    j h  h��h�!h�������ǅ����������T�������������  ��@���t!h8j h  h��j���������u̋����������������������������������������H��P���������������T�������P��h���P��d���Q��G���R��P���P������Q������R�H�P�l�Ѓ���������   t-��d��� u$��T�������P������R�T�P�l�Ѓ���G�����gu3��������   u%��T����j���P������P�P�Q�l�Ѓ����������-u!��������   ��������������������������P��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ��������   t ƅ����0��4�����Q������ǅ����   �*ǅ����   ��������   t��������   ������������% �  �#  ������ u�MQ��������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������l�����l��� u!hj h�  h��j�V�������u̃�l��� uI����    j h�  h��h�!h������ǅ����������T��������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�h���u!h�j h�  h��j�F�������u̃�h��� uI� ���    j h�  h��h�!h�������ǅ����������T����� ����������  �R  �1����������������d�����d���R��������x�����|�����
  ������%   �#  ������ u�MQ���������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������`�����`��� u!hj h�  h��j�"�������u̃�`��� uI�����    j h�  h��h�!h������ǅ����������T����������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�Q���������؉�\���u!h�j h�  h��j��������u̃�\��� uI�p����    j h�  h��h�!h��x�����ǅ����������T���������������  �  �1����������������X�����X���R���������x�����|�����  �������� �a  ��������@�'  ������ u�UR����������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������T�����T��� u!hj h�  h��j���������u̃�T��� uI�=����    j h�  h��h�!h�E�����ǅ����������T��������������  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������R��G���Pj��������������R����������؉�P���u!h�j h�  h��j���������u̃�P��� uI�-����    j h�  h��h�!h��5�����ǅ����������T��������������s  ��  �3����������������L�����L���P����������x�����|����&  ������ u!�MQ�^����������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������H�����H��� u!hj h�  h��j��������u̃�H��� uI�����    j h�  h��h�!h������ǅ����������T����g����������Z  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q�����������؉�D���u!h�j h�  h��j��������u̃�D��� uI�����    j h�  h��h�!h�������ǅ����������T����W����������J  �  �5����������������@�����@���R�]����������x�����|����V  ��������@�%  ������ u�MQ�$��������x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������<�����<��� u!hj h  h��j��������u̃�<��� uI������    j h  h��h�!h�������ǅ����������T����0����������#  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�8���u!h�j h  h��j�o�������u̃�8��� uI������    j h  h��h�!h��������ǅ|���������T���� �����|����
  �{  �2����������������4�����4���R�&��������x�����|����"  ������ u�EP�������3ɉ�x�����|�����  ������ |������d}ǅ����   �
ǅ����    ��������0�����0��� u!hj h0  h��j�Y�������u̃�0��� uI�����    j h0  h��h�!h������ǅx���������T����
�����x�����  ��@��� �
  �������������� uE��������Ǆ����   ����������G������������������������������   ������Q��G���Rj��������������Q����������؉�,���u!h�j h4  h��j�I�������u̃�,��� uI�����    j h4  h��h�!h�������ǅt���������T����������t�����  �U  �3����������������(�����(���R� �����3ɉ�x�����|�����������@tG��|��� >|	��x��� s3��x����؋�|����� �ى�p�����t�����������   ���������x�����p�����|�����t����������� �  u(������%   u��p�����t����� ��p�����t�����d��� }ǅd���   �%�����������������d���   ~
ǅd���   ��p����t���u
ǅ����    ��O�����������d�����d�������d�������p����t�����   �������RP��t���P��p���Q������0�������������RP��t���R��p���P�z�����p�����t���������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�s  ��l��� �B  ��������@t[��������   tƅ����-ǅ����   �:��������tƅ����+ǅ����   ���������tƅ���� ǅ����   ������+�����+�������$�����������u��L���Q�UR��$���Pj �m  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��$���Qj0�  �������� ��   ������ ��   ǅ���    �������� �����������������������������������   �� ���f�f������������Rj�����P�����Q�n������������ ������� �������� u	����� uǅL��������-��|���P��L���Q�UR�����P�����Q�  ���S����(��|���R��L���P�MQ������R������P�P  ����L��� |'��������t��L���R�EP��$���Qj ��  �������� tj������R�O�����ǅ����    ������8��� t��8���tǅ����    �
ǅ����   ���������������� u!h�j h�  h��j��������u̃���� uI�����    j h�  h��h�!h�������ǅp���������T����a�����p����T  �������%  ��@��� �  ǅ����    ���������������������;�x�����  �����������������������������������������  �������$������������E�������MQ��������  ���������E�������MQ�k������_  ���������E�������MQ�������;  ���������E�������MQ�������  ���������E�������MQ�r�������   ���������E�������MQ�:�������   ���������E�������MQ��������h�����l����   3�tǅ����   �
ǅ����    ���������������� u!hpj h.	  h��j��������u̃���� uF������    j h.	  h��h�!hp�������ǅd���������T����1�����d����'������s�����L�����`�����T���������`����M�3�������]Ë�����������P���r���a�P����� �I ���������� �����|�����������e������!���   	
�������2�V���z��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�������E��}��u�M�������U����M���]����������������������������������������������̋�U��E�M���M��~!�UR�EP�MQ�	������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��w�U�    �E�M���M��~N�U��E��MQ�UR�E�P�z������M���M�U�:�u�E�8*u�MQ�URj?�O�������뢋E�8 u�M�U����]��������������������������������������������������̋�U��E����U�
�E��A��Q�]�����������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �j����E�    �EP�Y   ���E��E������   ��G���ËE�M�d�    Y_^[��]������������������������������������������̋�U����\�P�l�E��X�Q�l�E��U�;U�r�E�+E�����s3���   j�M�Q�������E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r"j}h�!j�E�P�M�Q�W������E��}� u:�U���U�E�;E�r%h�   h�!j�M�Q�U�R�!������E��}� u3��Q�E�+E����M����U��E��E��M�Q���\��UR���M���U����U��E�P���X��E��]�����������������������������������������������������������������������������������������������̋�U��EP�^���������؃�]��������������������̋�U��Qh�   h�!jjj �������E��E�P���\��\��X��}� u�   ��U��    3���]������������������������̋�U��j���������tj���������u#�=��uh�   �������h�   ������]�������������������������̋�U��Q�E�    �	�E����E��}�s�M��U;�H,u�E���L,���3���]�������������������������������̋�U���   ���3ŉE�EP�������E��}� ��  �E�    �}�   tN�}�   tE�}t?�M�Qj j j j������������������ t������t���E�   ��E�   �}� ��  j��������tj����������   �=����   j����E�}� tq�}��tk�E�    �	�U���U�}��  s%�E�M�U��J�������U�E��P��u����E� j �U�R������P�A�����P������Q�U�R�@��  �}�   ��  ǅ������������-x����  +ȉ�����������������j h  h1h�0h 0h�/h  hx��������P�x�����3�������f��  h  ������Rj ����u:j h  h1h�0hH/hT�������P������Q������P������������R�����������<vk������P��������������TA�������j h  h1h�0h�.jh�������+�������������+�Q������R�������P������j h  h1h�0h.h�h  hx��M�����P�_�����j h  h1h�0hx-�E�Ph  hx�������P�*�����h  h -hx��d������M�3��߷����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��h�������]���������̋�U��j�hبh9�d�    P���SVW���1E�3�P�E�d�    �e��Y����@x�E�}� t#�E�    �U��E�������   Ëe��E����������M�d�    Y_^[��]��������������������������������̋�U��Q������@|�E��}� t�U��ڽ����]�������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �e���P�l�E�}� t#�E�    �U��E�������   Ëe��E������W����M�d�    Y_^[��]��������������������������������������������̋�U��E���]�����������������̋�U���$V���P�l�E�3Ƀ} ���M��}� uh�2j jDhH2j�b�������u̃}� u0������    j jDhH2h42h�2��������   �  �E�     �}� �_  h2� �E�}� ut3�t	�E�   ��E�    �U��U�}� uh�1j jPhH2j�ǹ������u̃}� u0�(����    j jPhH2h42h�1�3������   ��   h�1�M�Q�T�E��}� ��   3�t	�E�   ��E�    �E܉E�}� uh�1j jVhH2j�7�������u̃}� uD��P�F������������0j jVhH2h42h�1��������P�������V�U�R���E�膾���E��E�Ph����;E�t
�M�Q��j�UR�U���u�����    �	���� �3�^��]����������������������������������������������������������������������������������������������������������������������������������������̋�U���   ���3ŉE�}��  �E�E���p����M�ǅd���    ǅh����   ��h���R�E�P�MQ�UR�EP�S�������l�����l��� ��   ����zt�  j j �MQ�UR�EP��������h�����h��� u��   j^h4jj��h���Q��������E��}� u��   ǅd���   ��h���R�E�P�MQ�UR�EP賱������l�����l��� u�   jih4jj��l���Q�}������U���E��8 u�]j jlh�3ht3h�2��l�����Q�U�R��l���P�M��R�V�����P�Y�������d��� tj�E�P������3��-  ��d��� tj�M�Q����������  �  �}��   �U��\�����\����     j j �MQ�UR����`�����`��� u�Zh�   h4jj��`���P��������\������\����: u�(��`���P��\����R�EP�MQ����u�3��mj��\����P���������\����    ����I�D�} u>ǅX���    j��X���R�E    P�MQ����u�����U��X����3������M�3��گ����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E���]�����������������̋�U��jj �EP�MQ��  ��]���������������������̋�U��jj �EPj ��  ��]�������̋�U��jj �EP�MQ�  ��]���������������������̋�U��jj �EPj �|  ��]�������̋�U��jj �EP�MQ�Z  ��]���������������������̋�U��jj �EPj �,  ��]�������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj ��  ��]��������������������̋�U��jh  �EP�MQ�  ��]������������������̋�U��jh  �EPj �y  ��]��������������������̋�U��jh  �EP�MQ�G  ��]������������������̋�U��jh  �EPj �  ��]��������������������̋�U��jhW  �EP�MQ��  ��]������������������̋�U��jhW  �EPj �  ��]��������������������̋�U��jj�EP�MQ�  ��]���������������������̋�U��jj�EPj �\  ��]�������̋�U��jj �EP�MQ�:  ��]���������������������̋�U��jj �EPj �  ��]�������̋�U��jj �EP�MQ��   ��]���������������������̋�U��jj �EPj �   ��]�������̋�U����EP�M�迺���M��I����x t8�M��;����H�y�  u$jj �UR�EP�i   ���E�M������E���E�    �M������E��]��������������������������������̋�U��j �EP�f�����]�����������̋�U��j�h�.d�    P�����3�P�E�d�    �EP�M������E�    �M�M�M��l����P�E�L#Mu;�} t�M��N�������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M������E��M�d�    Y��]��������������������������������������������������������������̋�U��E�U��DV�u�     j�E�P3�NVf�
����u3�^��]ËM�U�E�QRP����t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D$+�3�3ۅ�t�;�r	��+�;p�rC��(;�r�;�t[C�=�� u �=�� uH�  �����t:�������h�4P�T3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�RhP�V�Ѕ��p  �M��R VVV�E�PWS�҅��K  �M�u���@h�U�R�Є��(  �M�;��  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�wE�;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj ��P�T�����   �M���RV�E�Pj j j �E�P�҄�tR+}�;>rK�M��   ;�v
;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj ��P�d�M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  ���3ŉE��=�� t3��M�3��R�����]������   ����   VWhp4���= �5���t?h  ������QP�օ�t,h  ������R������P��  ����t������Q�ׅ�uBh  ������Rj �օ�t,h  ������P������Q�  ����t������R�ׅ�u3�_^�M�3�营����]����������������������������������������������������������������̋�U���  ���3ŉE�Vh2� ����u^�M�3�������]�W�=Tht5V�׉�������u_^�M�3�������]�Sh`5V�׋؅�t4hP5V�׋���t&������Pjj h�4h  ���������tV��[_3�^�M�3�蛤����]Í�����Q������������R������Pj h�4Qǅ����  �Ӌ�����R����V����u�������u��������u����r�Hf9�E����u�f��E����\t�\   f��E����@���+Ѓ��\����H��  �M����T4�X4��E������\4�H�`4�P�d4�H�h4�Pf�l4�Hf�P������P� �M�[_3�^薣����]����������������������������������������������������������������������������������������������������������������������̋�U���  ���3ŉE��EV�uh   ������Qh   ������Rh   ������Qj�U�RP�ҥ����$��t3�^�M�3�輢����]�h�5������j	P�7�������u�h�5������jQ��������u�������R������P�E������Q�U�RPV�0����M������3�@^�N�����]��������������������������������������������������������������̋�U����E%�����E�M#M��������   �} tj j �ɦ�����U�3�t	�E�   ��E�    �M��M��}� uhX6j j1h�5j��������u̃}� u-�Q����    j j1h�5h�5hX6�\������   �/�} t�EP�MQ�=������U���EP�MQ�&�����3���]����������������������������������������������������������������̋�U����EP�M������M�虥����t2�M�荥������   ~�M��z���Ph  �UR��������E��h  �EP�M��R���P謟�����E�M�M�M��Ž���E��]��������������������������������������������̋�U��=�� uh  �EP��������j �MQ誳����]�������������̋�U����EP�M������M�詤����t/�M�蝤������   ~�M�芤��Pj�UR�������E��j�EP�M��h���P������E�M�M�M��ۼ���E��]����������������������������������̋�U��=�� uj�EP�(�������j �MQ�f�����]����������������̋�U����EP�M��?����M��ɣ����t/�M�轣������   ~�M�誣��Pj�UR�0������E��j�EP�M�舣��P�������E�M�M�M�������E��]����������������������������������̋�U��=�� uj�EP�H�������j �MQ�6�����]����������������̋�U����EP�M��_����M�������t/�M��ݢ������   ~�M��ʢ��Pj�UR�P������E��j�EP�M�訢��P�������E�M�M�M������E��]����������������������������������̋�U��=�� uj�EP�h�������j �MQ�w�����]����������������̋�U����EP�M������M��	�����t2�M����������   ~�M�����Ph�   �UR�m������E��h�   �EP�M��¡��P�������E�M�M�M��5����E��]��������������������������������������������̋�U��=�� uh�   �EP�u�������j �MQ�5�����]�������������̋�U����EP�M�菫���M�������t/�M���������   ~�M������Pj�UR耴�����E��j�EP�M��ؠ��P�2������E�M�M�M��K����E��]����������������������������������̋�U��=�� uj�EP蘝������j �MQ诜����]����������������̋�U����EP�M�诪���M��9�����t/�M��-�������   ~�M�����Pj�UR蠳�����E��j�EP�M������P�R������E�M�M�M��k����E��]����������������������������������̋�U��=�� uj�EP踜������j �MQ�������]����������������̋�U����EP�M��ϩ���M��Y�����t2�M��M�������   ~�M��:���Ph  �UR轲�����E��h  �EP�M�����P�l������E�M�M�M�腷���E��]��������������������������������������������̋�U��=�� uh  �EP�ś������j �MQ������]�������������̋�U����EP�M��ߨ���M��i�����t2�M��]�������   ~�M��J���PhW  �UR�ͱ�����E��hW  �EP�M��"���P�|������E�M�M�M�蕶���E��]��������������������������������������������̋�U��=�� uhW  �EP�՚������j �MQ������]�������������̋�U����EP�M������M��y�����t2�M��m�������   ~�M��Z���Ph  �UR�ݰ�����E��h  �EP�M��2���P茗�����E�M�M�M�襵���E��]��������������������������������������������̋�U��=�� uh  �EP��������j �MQ������]�������������̋�U����EP�M�������M�艜����t/�M��}�������   ~�M��j���Pj �UR�������E��j �EP�M��H���P袖�����E�M�M�M�軴���E��]����������������������������������̋�U��=�� uj �EP��������j �MQ賮����]����������������̋�U��}�   ���]��������������̋�U��E��]���̋�U��Q�EP�MQ�U�������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP�Z�������u�}_t	�E�    ��E�   �E���]�������������̋�U��Q�EP�MQ�z�������u�}_t	�E�    ��E�   �E���]�������������������������̋�U��Q�EP诚������u�M��_t	�E�    ��E�   �E���]�������������������������̋�U��E�� ]���̋�U���4�EP�M�诤���}   ��   �M��,�����t/�M�� �������   ~�M�����Pj�UR蓭�����E��j�EP�M�����P�E������Ẽ}� t,�M��љ������   �E��M��M��D����E��*  ��U�U܍M��,����E��  �M�菙��� ���   ~D�M��|���P�M�����   Q�D�������t"�U�����   �U��E�E��E� �E�   ��<���� *   �M�M��E� �E�   j�M�������BPj�M�Q�U�R�E�Ph   �M��������QR�M�����P账����$�E�}� u�E�E؍M��X����E��A�}�u�M��MԍM��>����E��'��U��E���ЉUЍM������E���M�������]����������������������������������������������������������������������������������������������������������������������������̋�U��Q�=�� u$�}A|�}Z�E�� �E���M�M��E���j �UR�j�������]���������������������������̋�U���@���3ŉE��E�    �E�    �EP�M������M��q���Pj j j j �MQ�U�R�E�P������ �E��MQ�U�R�g������E��E���u8�}�u�E�   �M�讯���E��j��}�u�E�   �M�蒯���E��N�:�M���t�E�   �M��t����E��0��U���t�E�   �M��V����E���E�    �M��B����E��M�3��ߑ����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�ř����]�������̋�U���@���3ŉE��E�    �E�    �EP�M��w����M�����Pj j j j�MQ�U�R�E�P譧���� �E��MQ�U�R�������E��E���u8�}�u�E�   �M��>����E��j��}�u�E�   �M��"����E��N�:�M���t�E�   �M������E��0��U���t�E�   �M������E���E�    �M��ҭ���E��M�3��o�����]�������������������������������������������������������������������������������̋�U��j �EP�MQ�i�����]�������̋�U���@���3ŉE��E�    �E�    �EP�M������M�葔��Pj j j j �MQ�U�R�E�P�=����� �E��MQ�U�R読�����E��E���u8�}�u�E�   �M��ά���E��j��}�u�E�   �M�責���E��N�:�M���t�E�   �M�蔬���E��0��U���t�E�   �M��v����E���E�    �M��b����E��M�3��������]�������������������������������������������������������������������������������̋�U��j �EP�MQ������]�������̋�U����E�E��M�Q�U�3��} ���E�}� uhl�j j7hX7j裓������u̃}� u0�����    j j7hX7h<7hl��������   �$  3�;U��؉E�uh��j j8hX7j�A�������u̃}� u0袪���    j j8hX7h<7h��譤�����   ��  �U� 3��} ����#E��;E��ىM�uh�6j j=hX7j�ɒ������u̃}� u0�*���� "   j j=hX7h<7h�6�5������"   �J  3��} ���E�}� uh�6j j>hX7j�c�������u̃}� u0�ĩ���    j j>hX7h<7h�6�ϣ�����   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R�m�������P�E��P�MQ������3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���,���3ŉE��EP�M�Q还�����U�Rj j���ċMԉ�U؉Pf�M�f�H�j������U�B�E�M��U��E�Pj j(hX8h<8h�7�M�Q�UR�EP蒨����P�Ӛ�����M�U�Q�E�M�3�蓊����]���������������������������������������������������̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]���������������������������������������������������������������������������������������������̋�U�������E��M�����Ƀ��M�uh�9j j*h9j�ʍ������u̃}� u+�+����    j j*h9h�8h�9�6������E���E����E���]��������������������������������̋�U����]����̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3������������������̋�U��j�^�����]���������������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ����������������������������XY�$�����������XY�$�����������XY�$����������̋�U���SVWd�5    �u��E�O;j �EP�M�Q�UR�g����E�H����U�Jd�=    �]��;d�    _^[��]� ����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�%����� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�՝���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ腝���� �E�_^[�E���]��������������������̋�U��E�HQ�U�B(Pj �M�QR薍����]� �����������������������̋�U����E�    �E�P=����M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ�D����E�E�d�    �E��]����������������������������������̋�U��Q��E�H3M跄��j �MQ�U�BP�M�QRj �EP�M�QR�EP�R����� �E��E���]��������������������̋�U���8S�}#  u�n>�M��   ��   �E�    �E��>����M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M��u������   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]��������������������������������������������������������������������̋�U��QS��E�H3M�&����M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ蠚���� �U�z$ u�EP�MQ诚��j j j j j �U�Rh#  �u������E��]�c�k ��   [��]���������������������������������������������������̋�U��Q�} �E�HSV�pW�M�����|8����u�0����E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v�����M�_��^��[��]��������������������������������̋�U��EV�u��P������   �N�B������   ��^]��������������������̋�U���������   ��t�M9t�@��u��   ]�3�]�������������������̋�U��V�؎���u;��   u�Ȏ���N���   ^]�跎�����   �x t�H;�t���x u�^]�����V�P^]�������������������������̋�U����EP�M������M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M��Y���P�.   ��$�E�M��ҝ���E��]�������������������������̋�U��� �} ~,�EP�MQ�%  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R��E��}� u3���  �}� ~63�u2�����3��u���r#h��  �M��T	R������P�,������E���E�    �E�E�}� u3��  �M�Q�U�R�EP�MQj�U$R���u
�Y  �T  j j �E�P�M�Q�UR�EP���E��}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR����u
��   ��   ��   �E��E�}� ~63�u2�����3��u��r#h��  �U�DP�������P�%������E���E�    �M��M��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ����u�V�T�}  u+j j j j �U�R�E�Pj �M$Q���E��}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P���E��}� t�M�Q�D������U�R�8������E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U����EP�M��ߋ���M$Q�U R�EP�MQ�UR�EP�MQ�M��M���P�2   �� �E�M��ƙ���E��]�����������������������������̋�U����E�    �} u�E��Q�Uj j �EP�MQ3҃}$ ��   R�EP��E�}� u3��   3�u2�}� ~,�}����w#h��  �U�DP�;�����P�b������E���E�    �M�M��}� u3��a�U���Rj �E�P�x������M�Q�U�R�EP�MQj�UR��E��}� t�EP�M�Q�U�R�EP���E��M�Q诖�����E���]�����������������������������������������������������������������������̋�U��Q�E�x  toj?h�:jhd  j�Ֆ�����E��}� u
�   �   �MQ�U�R��   ����t!�E�P�M�����j�M�Q�$������   �}�U�ǂ�      ��E����E���   ��tJ�M���   �´   R����u0�E���   ���    hp:j jOh�9j�|������u̋E�M����   3���]����������������������������������������������������������������̋�U����E�    �E�HB�M��U�BD�E��} u�����  �M�M��E�    �U��Rj1�E�Pj�M�Q詂����E�E�U��Rj2�E�Pj�M�Q舂����E�E�U��Rj3�E�Pj�M�Q�g�����E�E�U��Rj4�E�Pj�M�Q�F�����E�E�U��Rj5�E�Pj�M�Q�%�����E�E�U��Rj6�E�Pj�M�Q������E�E�URj7�E�Pj�M�Q������E�E�U�� Rj*�E�Pj�M�Q�Ł����E�E�U��$Rj+�E�Pj�M�Q褁����E�E�U��(Rj,�E�Pj�M�Q胁����E�E�U��,Rj-�E�Pj�M�Q�b�����E�E�U��0Rj.�E�Pj�M�Q�A�����E�E�U��4Rj/�E�Pj�M�Q� �����E�E�U��Rj0�E�Pj�M�Q�������E�E�U��8RjD�E�Pj�M�Q�ހ����E�E�U��<RjE�E�Pj�M�Q轀����E�E�U��@RjF�E�Pj�M�Q蜀����E�E�U��DRjG�E�Pj�M�Q�{�����E�E�U��HRjH�E�Pj�M�Q�Z�����E�E�U��LRjI�E�Pj�M�Q�9�����E�E�U��PRjJ�E�Pj�M�Q������E�E�U��TRjK�E�Pj�M�Q������E�E�U��XRjL�E�Pj�M�Q������E�E�U��\RjM�E�Pj�M�Q�����E�E�U��`RjN�E�Pj�M�Q�����E�E�U��dRjO�E�Pj�M�Q�s����E�E�U��hRj8�E�Pj�M�Q�R����E�E�U��lRj9�E�Pj�M�Q�1����E�E�U��pRj:�E�Pj�M�Q�����E�E�U��tRj;�E�Pj�M�Q��~����E�E�U��xRj<�E�Pj�M�Q��~����E�E�U��|Rj=�E�Pj�M�Q�~����E�E�U�   Rj>�E�Pj�M�Q�~����E�E�U�   Rj?�E�Pj�M�Q�e~����E�E�U�   Rj@�E�Pj�M�Q�A~����E�E�U�   RjA�E�Pj�M�Q�~����E�E�U�   RjB�E�Pj�M�Q��}����E�E�U�   RjC�E�Pj�M�Q��}����E�E�U�   Rj(�E�Pj�M�Q�}����E�E�U�   Rj)�E�Pj�M�Q�}����E�E�U�    Rj�E�Pj�M�Q�i}����E�E�U�¤   Rj �E�Pj�M�Q�E}����E�E�U�¨   Rh  �E�Pj�M�Q�}����E�E�U�°   Rh	  �E�Pj �M�Q��|����E�E�U�E����   �M���   Qj1�U�Rj�E�P��|����E�E�M���   Qj2�U�Rj�E�P�|����E�E�M���   Qj3�U�Rj�E�P�|����E�E�M���   Qj4�U�Rj�E�P�[|����E�E�M���   Qj5�U�Rj�E�P�7|����E�E�M���   Qj6�U�Rj�E�P�|����E�E�M���   Qj7�U�Rj�E�P��{����E�E�M���   Qj*�U�Rj�E�P��{����E�E�M���   Qj+�U�Rj�E�P�{����E�E�M���   Qj,�U�Rj�E�P�{����E�E�M���   Qj-�U�Rj�E�P�_{����E�E�M���   Qj.�U�Rj�E�P�;{����E�E�M���   Qj/�U�Rj�E�P�{����E�E�M���   Qj0�U�Rj�E�P��z����E�E�M���   QjD�U�Rj�E�P��z����E�E�M���   QjE�U�Rj�E�P�z����E�E�M���   QjF�U�Rj�E�P�z����E�E�M���   QjG�U�Rj�E�P�cz����E�E�M��   QjH�U�Rj�E�P�?z����E�E�M��  QjI�U�Rj�E�P�z����E�E�M��  QjJ�U�Rj�E�P��y����E�E�M��  QjK�U�Rj�E�P��y����E�E�M��  QjL�U�Rj�E�P�y����E�E�M��  QjM�U�Rj�E�P�y����E�E�M��  QjN�U�Rj�E�P�gy����E�E�M��  QjO�U�Rj�E�P�Cy����E�E�M��   Qj8�U�Rj�E�P�y����E�E�M��$  Qj9�U�Rj�E�P��x����E�E�M��(  Qj:�U�Rj�E�P��x����E�E�M��,  Qj;�U�Rj�E�P�x����E�E�M��0  Qj<�U�Rj�E�P�x����E�E�M��4  Qj=�U�Rj�E�P�kx����E�E�M��8  Qj>�U�Rj�E�P�Gx����E�E�M��<  Qj?�U�Rj�E�P�#x����E�E�M��@  Qj@�U�Rj�E�P��w����E�E�M��D  QjA�U�Rj�E�P��w����E�E�M��H  QjB�U�Rj�E�P�w����E�E�M��L  QjC�U�Rj�E�P�w����E�E�M��P  Qj(�U�Rj�E�P�ow����E�E�M��T  Qj)�U�Rj�E�P�Kw����E�E�M��X  Qj�U�Rj�E�P�'w����E�E�M��\  Qj �U�Rj�E�P�w����E�E�M��`  Qh  �U�Rj�E�P��v����E�E�E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��} u�W  j�E�HQ��}����j�U�BP��}����j�M�QR��}����j�E�HQ��}����j�U�BP�}����j�M�QR�}����j�E�Q�}����j�U�B P�}����j�M�Q$R�t}����j�E�H(Q�c}����j�U�B,P�R}����j�M�Q0R�A}����j�E�H4Q�0}����j�U�BP�}����j�M�Q8R�}����j�E�H<Q��|����j�U�B@P��|����j�M�QDR��|����j�E�HHQ��|����j�U�BLP�|����j�M�QPR�|����j�E�HTQ�|����j�U�BXP�|����j�M�Q\R�u|����j�E�H`Q�d|����j�U�BdP�S|����j�M�QhR�B|����j�E�HlQ�1|����j�U�BpP� |����j�M�QtR�|����j�E�HxQ��{����j�U�B|P��{����j�M���   R��{����j�E���   Q��{����j�U���   P�{����j�M���   R�{����j�E���   Q�{����j�U���   P�u{����j�M���   R�a{����j�E���   Q�M{����j�U���   P�9{����j�M���   R�%{����j�E���   Q�{����j�U���   P��z����j�M���   R��z����j�E���   Q��z����j�U���   P��z����j�M���   R�z����j�E���   Q�z����j�U���   P�z����j�M���   R�qz����j�E���   Q�]z����j�U���   P�Iz����j�M���   R�5z����j�E���   Q�!z����j�U���   P�z����j�M���   R��y����j�E���   Q��y����j�U���   P��y����j�M���   R�y����j�E���   Q�y����j�U��   P�y����j�M��  R�y����j�E��  Q�my����j�U��  P�Yy����j�M��  R�Ey����j�E��  Q�1y����j�U��  P�y����j�M��  R�	y����j�E��   Q��x����j�U��$  P��x����j�M��(  R��x����j�E��,  Q�x����j�U��0  P�x����j�M��4  R�x����j�E��8  Q�}x����j�U��<  P�ix����j�M��@  R�Ux����j�E��D  Q�Ax����j�U��H  P�-x����j�M��L  R�x����j�E��P  Q�x����j�U��T  P��w����j�M��X  R��w����j�E��\  Q��w����j�U��`  P�w����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���VW�E�    �E�    �E�E��E�    �M�y u�U�z �  jeh�;jjPj�,~�����E�}� u
�   ��  �E���   �   �}��jqh�;jj�8a�����E�}� uj�M�Q�lu�����   �z  �U��    �E�x �:  j}h�;jj��`�����E��}� u&j�M�Q�"u����j�U�R�u�����   �"  �E��     �M�Q>�U��E�Pj�M�Qj�U�R�j����E�E�E��Pj�M�Qj�U�R�dj����E�E�E��Pj�M�Qj�U�R�Cj����E�E�E��0Pj�M�Qj�U�R�"j����E�E�E��4Pj�M�Qj�U�R�j����E�E�t0�E�P�fx����j�M�Q�9t����j�U�R�+t��������;  �E�HQ�  ���@�E�    �U�8���M�<��Q�E�@��H�U�h��B0�M�l��Q4�E��    �}� t	�M��   ��E�    �E�    �E�8��U���    tA�E���   Q����u-�U���    w!hx;j h�   h ;j�$e������u̋M���    t<�U���   P����u(j�M���   R�"s����j�E���   Q�s�����U�E����   �M�U쉑�   �E�M䉈�   3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�   �E�;8�tj�U�P�?q�����M�Q;<�tj�E�HQ� q�����U�B;@�tj�M�QR�q�����E�H0;h�tj�U�B0P��p�����M�Q4;l�tj�E�H4Q��p����]�����������������������������������������������������̋�U���VW�E�    �E�E��E�    �M�y u�U�z �W  jSh�<jjPj�x�����E�}� u
�   ��  jYh�<jj��[�����E��}� uj�E�P�p�����   ��  �M��    �U�z �d  jeh�<jj�[�����E�}� u&j�E�P�o����j�M�Q�o�����   �s  �U��    �E�H8�M��E�    �U��Rj�E�Pj�M�Q�e����E�E�U��Rj�E�Pj�M�Q��d����E�E�U��Rj�E�Pj�M�Q��d����E�E�U��Rj�E�Pj�M�Q�d����E�E�U��Rj�E�Pj�M�Q�d����E�E�U�� RjP�E�Pj�M�Q�pd����E�E�U��$RjQ�E�Pj�M�Q�Od����E�E�U��(Rj�E�Pj �M�Q�.d����E�E�U��)Rj�E�Pj �M�Q�d����E�E�U��*RjT�E�Pj �M�Q��c����E�E�U��+RjU�E�Pj �M�Q��c����E�E�U��,RjV�E�Pj �M�Q�c����E�E�U��-RjW�E�Pj �M�Q�c����E�E�U��.RjR�E�Pj �M�Q�hc����E�E�U��/RjS�E�Pj �M�Q�Gc����E�E�U��8Rj�E�Pj�M�Q�&c����E�E�U��<Rj�E�Pj�M�Q�c����E�E�U��@Rj�E�Pj�M�Q��b����E�E�U��DRj�E�Pj�M�Q��b����E�E�U��HRjP�E�Pj�M�Q�b����E�E�U��LRjQ�E�Pj�M�Q�b����E�E�t@�U�R�q����j�E�P�l����j�M�Q�l����j�U�R�l�����   �b  �E�HQ�  ����   �8��}��U���   �M���E���   �U�A�B�M���   �E�J�H�U���   �M�P0�Q0�E���   �U�A4�B4�M��   �}� t	�U��   ��E�    �E�    �E�8��E���    tA�M���   R����u-�E���    w!hx<j h�   h <j�m]������u̋U���    t<�E���   Q����u(j�U���   P�kk����j�M���   R�Wk�����E�M䉈�   �U�E����   �M�U艑�   3�_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]���������������������������������̋�U��} u�  �E�H;D�tj�U�BP��h�����M�Q;H�tj�E�HQ��h�����U�B;L�tj�M�QR�h�����E�H;P�tj�U�BP�h�����M�Q;T�tj�E�HQ�h�����U�B ;X�tj�M�Q R�bh�����E�H$;\�tj�U�B$P�Ch�����M�Q8;p�tj�E�H8Q�$h�����U�B<;t�tj�M�Q<R�h�����E�H@;x�tj�U�B@P��g�����M�QD;|�tj�E�HDQ��g�����U�BH;��tj�M�QHR�g�����E�HL;��tj�U�BLP�g����]�����������������������������������������������������������������������������������������������������������̋�U����&a���E��E��Hl�M��U�;D�t�E��Hp#��u�g���E������]�����������������������������̋�U�졤�]����̋�U����`���E��E��Hl�M��U�;D�t�E��Hp#��u�&g���E��U����   ��]�������������������������̋�U���EP�MQ�b����]�������̋�U��Q�E=��  u3��G�M��   }�U����P�M#��&�U�Rj�EPj����u3�f�M��E��U#�]��������������������������������̋�U���EP�MQ��a����]�������̋�U��j
j �EP�Z����]���������̋�U��EPj
j �MQ��[����]���������������������̋�U��EP��m����]�������������̋�U��EP�MQ�\����]���������̋�U��j
j �EP��U����]���������̋�U��EPj
j �MQ�h����]���������������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh�j jh�Fj�V������u̃}� u0�tm���    j jh�Fh�Fh��g�����   �J  �} u\�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U�E�Ph�   �M��Q�V����3���  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�U����3҃} �U��}� uhL�j jh�Fj��T������u̃}� u0�Ml���    j jh�Fh�FhL��Xf�����   �#  �M�M��U�U��}�u5�E��M���E���U����U��E���E��t�M����M�t���y�_����t&�U;Urh�j j+h�Fj�@T������u̋M��U���M���E����E��M���M��t�U����U�t�E���Et�} u�M�� �}� ��   �}�u�UU�B� �P   �?  �E�  �}�tI�}���t@�}v:�M��9��s����U��	�E���E܋M�Qh�   �U��R�T��������t3�t	�E�   ��E�    �U؉U�}� uh��j j>h�Fj�6S������u̃}� u-�j��� "   j j>h�Fh�Fh���d�����"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9��s����M���U+U����E+EԋM�Qh�   �U+U��E�LQ�S����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�hH�h9�d�    P���SVW���1E�3�P�E�d�    3��} ���E��}� uh$Hj jNh�Gj�(Q������u̃}� u-�h���    j jNh�Gh�Gh$H�b����3��   h�  �UR�ia����=�  ��؉E�uh@Gj jOh�Gj�P������u̃}� u*�h���    j jOh�Gh�Gh@G�$b����3��<j�Q�����E�    �UR�M�����E��E������   �j��]����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U�������E��=H� u3���   �}� u"�= � t��H����t3���   ����M��}� ��   �} ��   �UR�}R�����E��E��8 ��   �M��R�`R����;E�v{�E���U����=uj�M�Q�UR�E��Q�^������uPh�  �U���M��TR�_����=�  r!hPHj h�   h�Gj��N������u̋M���E��D��M����M��X���3���]�����������������������������������������������������������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    j�ZO�����E�    �EP�MQ�UR�EP�X   ���E��E������   �j�[����ËE�M�d�    Y_^[��]������������������������������������̋�U���3��} ���E��}� u!hJj h�   h�Gj�M������u̃}� u3��d���    j h�   h�Gh�IhJ��^�����   �   �U�    �} t�} w�} u�} t	�E�    ��E�   �E��E�}� u!h(Ij h�   h�Gj��L������u̃}� u3�Yd���    j h�   h�Gh�Ih(I�a^�����   �   �} t�U� �EP�@I�����E��}� u3��d�M�Q�O�������U��} u3��F�E�;Mv�"   �5j h�   h�Gh�Ih�H�U�R�EP�MQ��d����P�W����3���]��������������������������������������������������������������������������������������������������������̋�U��j j j�EP�MQ�UR��^����]���������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    j�zL�����E�    �EP�MQ�UR�EP�MQ�UR�`   ���E��E������   �j�X����ËE�M�d�    Y_^[��]��������������������������������������������̋�U���3��} ���E�}� u!h�Jj hX  h�Gj�J������u̃}� u3� b���    j hX  h�Gh�Jh�J�\�����   �2  �U�    �} t	�E�     3Ƀ} ���M��}� u!h�Jj h^  h�Gj�J������u̃}� u3�|a���    j h^  h�Gh�Jh�J�[�����   �   �EP�oF�����E��}� u3��   �M�Q��L�������E��UR�EP�MQj�U�R�<`�����M��U�: u��`���    ��`��� �Ej hr  h�Gh�Jh@J�E�P�M�Q�U�P��a����P�T�����} t�M�U��3���]����������������������������������������������������������������������������������������������������������������������̋�U���@���3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �M�y ��  �U�z u+�E��Ph  �M�Q0Rj �E�P�L������t�"  j^h�Kjj�B�����E�jbh�Kjjh�  �^�����E�jdh�Kjjh�  �^�����E�jfh�Kjjh�  �u^�����E�jhh�Kjjh  �Z^�����E�}� t�}� t�}� t�}� t�}� u�}  �M��    �U�U��E�    �	�E����E��}�   }�M��U���E����E��ۍM�Q�U�BP�0��u�&  �}�v�  �M܉Mă}�~S�U�U��	�E����E��M����t8�E��H��t-�U���E��	�M����M��U��B9E��M�M�� ���j j �U�BP�Ḿ�   Qh   �U�Rjj �S���� ��u�  j �E�HQh�   �Uȁ   Rh�   �E��Ph   �M�QRj �S����$��u�E  j �E�HQh�   �U��   Rh�   �E��Ph   �M�QRj �]S����$��u�  3��M�f���   �U��B �E��@ �M�Ɓ�    �U�Ƃ�    �}�~]�E�E��	�M����M��U����tB�M��Q��t7�E���M��	�U����U��E��H9M�� �  �E��M�f��A   ���h�   �Ú�   R�E�P��N����j�Mȁ�   Q�U�R�N����j�E�   P�M�Q�N�����U���    ��   �E���   Q������   3�uj j h�   h@Kj��D������u�j�M���   ���   R�
S����j�E���   ��   Q��R����j�U���   -�   P��R����j�M���   R��R�����E��    �M�UЉ��   �E�   �M���   �Ú��   �E���   �Mȁ��   �U���   �E��   �M���   �U�Eĉ��   j�M�Q�NR����3���   j�U�R�9R����j�E�P�+R����j�M�Q�R����j�U�R�R����j�E�P�R�����   �   �   �M���    tA�U���   P����u-�M���    w!h Kj h�   h@Kj�sC������u̋Eǀ�       �Mǁ�       � >�E���   ��B�U���   �D�M���   �Uǂ�      3��M�3��=����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�����I���E��E��Hl�M��U�;D�t�E��Hp#��u�FP���E��U����   ��]�������������������������̋�U��Q�} u
�V���E���E����   �U��E���]���������������������̋�U����6I���E��E��Hl�M��U�;D�t�E��Hp#��u�O���E��U��B��]����������������������������̋�U�����H���E��E��Hl�M��U�;D�t�E��Hp#��u�FO���E��U��B��]����������������������������̋�U����vH���E��E��Hl�M��U�;D�t�E��Hp#��u��N���E��E�����]����������������������������̋�U���]����̋�U���]����̋�U�����G���E��E��Hp����Ƀ��M��U�U��E����E��}�wC�M��$����U��Bp���M��Ap�   �U��Bp����M��Ap�   �   ��������u3�t	�E�   ��E�    �E�E�}� u!h�Mj h�   hhMj��>������u̃}� u.�_V���    j h�   hhMh8Mh�M�gP���������E���]Ð/�*��������������������������������������������������������������������������̋�U��j�h��h9�d�    P��SVW���1E�3�P�E�d�    �=D�@�tAj�>?�����E�    h@�hD���R�����D��E������   �j�K����ËM�d�    Y_^[��]�����������������������������������������������̋�U��j�hȩh9�d�    P��SVW���1E�3�P�E�d�    �} ��   j�>�����E�    �E�x t.�M�QR����u�E�x`�tj�M�QR�XK�����E������   �j�J����ËE�8 tcj�>�����E�   �M�R�P�����E�8 t#�M��: u�E�8@�t�M�R�8�����E������   �j�DJ����ËE� 𭺋M�A�j�UR�J�����M�d�    Y_^[��]�������������������������������������������������������������������������������������̋�U��EP�=����]�������������̋�U����E�    �} |�}�} u3��  he  hTNjjj�\R�����E��}� u�S���    3��  hj  hTNjjh�   �&R�����M���U��: u j�E�P�I������R���    3��8  hp  hTNjjh   ��Q�����E��M��U��Q�}� u0j�E��Q�LI����j�U�R�>I�����sR���    3���   h@��E��Q�P  ���UR�EP�M��R�z  ����u3�E��Q�nN�����U��P�6����j�M�Q��H�����E�    �x�U��BP�M���BP�%<������tDj�M��QR�H�����E��Q�N�����U��P�@6����j�M�Q�uH�����E�    ��U��B�    �M��Q�   �E���]���������������������������������������������������������������������������������������������������������������������������������̋�U��VW�} t0�} t*�E;Et"�u�6   �}�M�    �UR�XL����_^]�������������������������������̋�U��EP�MQ�_D����]���������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �E�    �%A���E�h�  hTNjjj�cO�����E�}� u�P���    3��   �G����I���E�M��Ql��E�M��Qh�Pj�9�����E�    �E�Q�aK�����E������   �j��E�����j�_9�����E�   �U�BP���E������   �j�E����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������̋�U����H��]����̋�U��j�h(�h9�d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �EԉE؃}� u!h�Nj h&  hhMj�!7������u̃}� u0�N���    j h&  hhMh�Nh�N�H����3��  �/?���E���E���U܋Bp���M܉Ap�E�    h1  hTNjjh�   �OM�����E�}� �  j�7�����E�   �U܋BlP�M�Q��������E�    �   �j�D����Ã}� ��   �UR�EP�M�Q��  ���E��}� ��   �} th���UR�c9������t
���   j�%7�����E�   �E�P�M܃�lQ�J�����U�R�I�����E܋Hp��u$�����u�E܋HlQhD��vJ�����
  �E�    �   �j�=C�������U�R�<I�����E�P�p1�����E������   ��M܋Qp���E܉PpËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��D����   ����D����   ����D����   ���]���������������������̋�U���   ���3ŉE��} tC�} t�EP�MQ�UR�  ����T�����E���M�TH��T�����T����E��|  ǅd���   ǅh���    �} �O  �M���L�'  �E�H��C�  �U�B��_�  �M��`���h�O��`���R�p,������\�����\��� t"��\���+�`�����X���t��\������;u3���  ǅl���   ���l�������l�����l���N��X���Q��`���R��l���k���HLQ�C������u"��l���k���HLP��5����9�X���u�뚋�\�������\���h�O��\���R�b+������X�����X��� u��\������;t3��$  ��l���|j h�  hhMh�OhO��X���R��\���Ph�   ��p���Q� 0����P�#=������X���Ƅp��� ��p���P��l���Q�UR��  ����t��h�������h�����\����X�����`�����`������t��`�������`�����`�������7�����h��� t�MQ��  ����P����
ǅP���    ��P����U��  �EPj j h�   ��p���Q�UR�E�����E��}� ��   ǅl���    ���l�������l�����l���|��l��� tn��l������U�D
HP��p���Q�p4������t;��p���R��l���P�MQ�  ����t��h�������h����
ǅd���    ���h�������h����l�����d��� t�MQ��  ���E��0��h��� t�UR�  ����L����
ǅL���    ��L����E���MQ�  ���E��E��M�3��+����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  ���3ŉE�ǅX���    ǅT���    �7����D�����D����  ��l���ǅH���   �MQ��@���R��L���Ph�   ��p���Q�UR�C������u3��  �E���M�THR��p���P�2������u�M���U�D
H�a  ��p���P�1��������T���h�  hTNj��T���Q�g(������X�����X��� u3��  �U���E�LH��8����U�E�L���<���j�Uk��E�L$Q��0���R�7�����E�H��\���j h  hhMhdPh�O��p���R��T�����P��X�����Q�eF����P�8������X������E���M�TH��L����E�M�T�j��L���R�Ek��M�T$R��6�����}�
  �E��@����H��H�����l����L���T����(�����,���ǅ`���    ���`�������`�����`���;�H�����   �U��`�����l����R;�uJ��`��� t=��`�����l������D���l�����A��`�����l�����(����Ћ�,����L��]�V��`�����l����ЋT���d�����h�����`�����l�����(�������,����T���d�����(�����h�����,����#�����`���;�H�����   j�E�HQ�U�BP��8���Qjh�Ljj �8���� ����   ǅ$���    ���$�������$�����$���s$��$�����E8������  ��$���f��U8�����h�   �(�P��8���Q�5������u��l����B   ���l����@    ���l����A    ��l����E�H�
�U��l����H���   �}u�U��@����B�MQ�Uk���PL�Ѓ���tG�M���U��8����D
Hj��X���Q�c9�����U�E��<����L��U��\����B3��   ��8�����t{�M���U�D
PP����uc3�uj j h[  hhMj��*������u�j�E���M�TPR��8����j�E���M�TTR��8�����E���M�DL    ��X��� t��X����   �E���M��X����TP�E���M�DH�M�3���$����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�    �E�    �E�    �E�U  ht  hTNj�E�P�"�����E�}� u3��  �M���M��U���U��E��  �M��   �E�   �	�U����U��E����M�THRh Q�E�k���HLQj�U�R�E�P�7!�����}�}kj h�  hhMh�Ph�Ph�O�M�Q�U�R�� ����P��2�����E������M�THR�E����M�THR�+������t�E�    �  �}� ��   �E�xP tD�M�QPR����u33�uj j h�  hhMj�'������u�j�U�BPP�5�����M�yT tD�U�BTP����u33�uj j h�  hhMj�7'������u�j�E�HTQ�X5�����U�BT    �E�@L    �M�U�QP�E�M��HH�E���   ��   j�U�R�5�����E�xP tD�M�QPR����u33�uj j h�  hhMj�&������u�j�U�BPP��4�����M�yT tD�U�BTP����u33�uj j h�  hhMj�\&������u�j�E�HTQ�}4�����U�BT    �E�@L    �M�AP    �U�BH    �E�@h�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����   ���3ŉE��y-���   �E�E��(�E��M�� �M�U��,�U��E�   �E��   �E��E��   �E�    �} u3��-  �} t�} u3��  �M���Cuv�E�H��ukj h�  hhMh\RhRhR�UR�EP�=����P�O/�����} t3ɋUf�
3��Mf�A3ҋEf�P�} t	�M�    �E�  �UR�K'�����E��}��   s0�EP�M�Q�f'�������  �UR�E�P�N'��������   ǅ@���    ǅD���    �MQ��H���R�I%������t3��  ��H���P�M�Q��H���R�P&������u3���   �E��H�U��
��H���P�M�Q�U�R�'�����E���t�}��   s�U��@����E���D����
ǅ@���k�j h�  hhMh\RhhQ��D�����Q��@���R�E�P�M�Q�� ����P��-�����} tj�U�R�EP�[,�����} tj�M�Q�UR�C,����j h  hhMh\RhQ�E�P�MQ�UR�A;����P�-�����E��M�3��K����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�]�������̋�U����E�E��E�    �	�M����M��U�;U}A�E����E�j h  hhMh4Th�R�M��Q�R�EP�MQ�B����P�O,������E�    ��]��������������������������������������������̋�U���h�   j �EP�!�����M���u3���  �E���.uX�U�B��tMj h*  hhMh0Xh0Wj�M��Qj�U�   R�����P�+�����Eƀ�    3��e  �E�    �	�M����M�h,W�UR�5�����E��}� u����1  �EE���M��}� uI�}�@sC�U���.t:j h8  hhMh0Xh8V�E�P�MQj@�UR������P��*�����   �}�uI�}�@sC�E���_t:j h;  hhMh0XhHU�M�Q�URj@�E��@P�����P�*�����_�}�uT�}�sN�M���t	�U���,u=j h>  hhMh0XhPT�E�P�MQj�U�   R�O����P�R*���������)�E���,u��M���u��U��E�L�M����3���]����������������������������������������������������������������������������������������������������������������������������������������̋�U��j hT  hhMh�XhXX�EP�MQ�UR�7����P�^)�����E�H@��t�U��@RhTXj�EP�MQ�e�����U���   ��t!�M���   QhPXj�UR�EP�6����]����������������������������������������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���������������������������̋�U��j�hh�h9�d�    P���SVW���1E�3�P�E�d�    �E������E������}�u!�#���     ��4��� 	   ��������  �} |�E;h�s	�E�   ��E�    �MԉM܃}� uh8�j jMhYj�������u̃}� u<� #���     �^4��� 	   j jMhYh Yh8��i.�����������C  �E���M���������D
������؉E�uh��j jNhYj�������u̃}� u<�"���     ��3��� 	   j jNhYh Yh����-�����������   �UR������E�    �E���M���������D
��t �MQ�UR�EP�MQ������E��U��F�Q3��� 	   ��!���     �E������E�����3�uh��j jYhYj�������u��E������   ��MQ������ËE��U�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��UR�$�����E�}��u;�2��� 	   3�u!h��j h�   hYj�������u̃������   �UR�E�P�M�Q�U�R���E��}��u#���E��}� t�E�P�[�����������>�M���U���������L����U���E���������L�E��U���]������������������������������������������������������������������������̋�U��j�h��h9�d�    P�ĘSVW���1E�3�P�E�d�    �} u3��   j�A������u3��oj�k�����E�    �EP�MQ� ��0/���URj �EP�MQ�UR�M��0���M��0���E� ��&���E������   �j�&����ËE�M�d�    Y_^[��]��������������������������������������������������������������̋�U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� �����������������̋�U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]�������������������̋�U��j�h��h9�d�    P�ĘSVW���1E�3�P�E�d�    �} u3��   j�������u3��pj������E�    �EP�MQ� ��p-���U R�EP�MQ�UR�EP�M��D.���M���.���E� ��M$���E������   �j��$����ËE�M�d�    Y_^[��]�������������������������������������������������������������̋�U��Q�M��M���-���M���,��-���E�$��$�� ��} t�U�,��E�(���(�    �,�    �M���,���U����E�0��M�4��8� �E���]� ��������������������������������������������̋�U���H�M��M��(���M�� ���=$� ��   �$����?uG�$��B��@u8� ���� ��U�R�����Ph�a�E�P�$����P�M�����v�$����?uS�$��H��$uEj �U�R�W'����P�M������M�������u�$�� ��M�Q�-����P�M������U�R�����P�M�����M������u	3��  �?�M��y����t�'����u� ����t�$�R�M��S����E�P�M��:���=(� u2�M��+�����,�jh ��,�Q�F!�����E��U��(��=(� ��   �,�P�(�Q�M���$���(��U�E�E�M����tY�E���� u0�U���U�E��  �M���M�U���� u�M���M�����U�E��
�U���U�E���E�띋M�U���(���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M�jPhH��M��#���H���]���������������̋�U���h�� ����tH�0�%�����0�j �M�Q������0���    �0��E�P�M�����E�  �  � ����?�t  � ���� �� ����?uK� ��H��?u=�U�R�o����� ����t� ���� ���E�P�M�L���E�9  �M�Q�\�����M�����E�M������E��M�������u�U�R�M�
���E��  � ������   � ����@��   �M�Q������M��$������   �8���tn�8� �E�P�M�Q�M����P�M����� ����@t>�M�Q�=����P�M���
���U�R�E�Ph�a�M�Q�M�������Y��P�M���
���)�U�R�E�Ph�a�M�Q�M��r�����.��P�M��
���}� t�M�����}� t�M��r���M��V����u�M��u����t�U�R�M�����E��   �   � ����t� ����@ut� ����t� ���� ��"����t:�}� u4�M��@����u(�M����P�M�Q��'�����U�R�M�e���E�U��E�P�MQ�'�����E�>�j�M����E�-�+� ����tj�M����E��j�M�z���E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U�� ����?uJ� ��B��$uj�MQ�� �����E�;�$� ���� �j j �EP��'�����E��j j�MQ�������E]�������������������������������̋�U���h���3ŉE� ����0�M�x5�}�	/� ���� ��E�P�MQ�������E�;  �6  �M��|��� ����?ubj �M�Q�" ����P�M����� ��� ���� ���@t)� ���� �� ������ك�Q�M�����  jh b� �R���  ����u�E� b� ���� ��9jh�a� �Q�ί  ����u�E��a� ���� ���E�    �}� ��   �E�P������.����twj�M�Q�M������U�R�,$����P�4����EЃ}� t�E�P�M�����:h�a�M����h�a�M�Q�U�R�E�P�M�Q���������"��P�M������:h�a�M��Q��h�a�U�R�E�P�M�Q�U�R�����������P�M�����N�E��t.� ����@u �M����P�M������ ���� ��j@h ��M�����P�M������M��t�������u�U�R���N���E�P�M����E�M�3�������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  �M��x���M��p���E�    �E�    � �������� ���� ����������������_�o  �������\��$�@�� ���� �j�M�7���E�  �M������M����   �U�R�;����Pj<�E�P�����P�M��
���M������ȃ�>u
j �M����j>�M�����} t�U�� ����u�U�R�M�C���E�  � ���� �� ��M�j j �U�R�����P�M�����Eܣ ��M��T����u*� ��Q���1u�E�Pj~�M�Q�\����P�M��J���M������u�U�R�M���	���E�P�M����E�v  �%  � ��Q���p_P�M��
���  �E�   � ��Q���T_P�M�������  � �������� ���� ����������������_��  ����������$���� ���� �j�M�b���E��  � ��B��� `Q�M��[���F  � ��B��� `Q�M�����E�  �  � ��B��� `Q�M�����M������U�R�M�z���E�F  ��  jhl^�E�P�7�����M��V���M�Q�M�F���E�  � ��B����_Q�M�J���E��  � ��B����_Q�M����j j �U�R�!����P�M��e���M��9����u�M��H
����tj�M�3���E�  �E�P�MQ�M�����E�{  �  �  � ��B����_Q�M��
��� ����uj�MQ�M�� ���E�4  � ����0�E�x�}�rj�M����E�  �M���xaR�M����� �������� ���� ������������������0�����������>  ������$�P�j �E�P� �����M�Q�UR�E�P��t���Qj ��|���R�M���������������E�^  �  �E�P�M�Q�M��x��j,��d���R��l���P��������7��P�M��h��j,��T���Q��\���R����������P�M��@��j,��D���P��L���Q�X����������P�M����j)��4���Rj ��<���P����������P�M�����j'�MQ�M�����E�  �;�U�R�EP�M�����E�w  �!� ���� �j�M�����E�T  ��  � ��B����_Q�M�������  � ���� ���� ���� ��� ��������������� t������0t!�N� ���� �j�M�s���E��  j hb�M�Q��������M������U�R�M�����E�  j�M�2���E�  �0  � ��������� ���� ���������������������A������������	��   ��������l��$�d�� ��Q���H`P�M�l����E�  � ��Q���H`P�M��J���� ����?u5��,���P�
����P�M����� ����@u� ���� ����$���Q������P�M�����hb�M��p���U�R�M����E��j�M����E�n�j�M�����E�]�j�M�����E�L�}� t
�M������-�M������u!�E�Ph@_�����Q�5����P�M������U�R�M�/���E��]ÍI ����Ƚ����� V�w�����	�'���I�ÿȿ������ 	

�����������'�        �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M������ ��� ���� ���@u� ��� ���� ���_tj�M����E�   � ���� �j �U�R������j �E�P������� ����t� ����@t� ���� ��ա ����u� ���� �j�M�*���E�� ���� ��M�Q�M�
���E��]��������������������������������������������������������������������̋�U����   �M��x���E� �M���������  � ������  � ����@��  �8���t�9���u�E�P�M��	���E�(  �M��2����uE�M�Qh�a�U�R�����P�M��4����E���t�M�Qj[�U�R�#����P�M������E� � ����?�  � ���� �� ����@�����@�����$��@�����@���%��  ��@��������$���� ��B��_ua� ��Q��?uR� ���� ��M�Q�U�Rj j �E�P������������P�M��\���� ����@u� ���� ��@�M�Q�U�Rj'�E�P�M�Q�����Pj`�U�R��������t���������P�M��������   � ���� ��M�Q�U�Rj j�E�P�S�������U���P�M��������   j@h ��M�����M�Qhb�U�R�����P�M�������������u�E�P��� ����w� ���� ��U�R��|���Pj]�M�Qj j�U�R������������������P�M��,����E��*�E�P��l���Q��t���R�@����������P�M�������.�E�P��\���Qj j��d���R�Z�������\���P�M����������� ����<�����<��� t��<���@tW�W�M��z����tj�M�������;�U�R��D���Ph�a��L���Qj��T����Z	�����'���������P�M��S�����
j�M������U�R�M����E��]Ð��!�2�n��� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���� ����uj�M�����E�T�R� ����?u3� ���� �j �U�R�����Pj-�EP� �����E��j �MQ�������E��]�������������������������������������̋�U���   V�E�    � ����Qu�E�8b� ���� �� ����uj�M����E�S  �N  � ����0��   � ����9��   �}� tG� �� ��/��E��U�� ���� ��U�R�E�P�M�����P�M�Q�U�R������E��4� �� ��/��E��U�� ���� ��U�R�E�P�M�����E��M��M�U�R�M�����E�  �  �E�    �E�    � ����@��   � ����uj�M�����E�L  �W� ����A|7� ����P*�E��U���;����ȋ� ����A���M��u��j�M����E��   � ���� ��e���� ��� ���� ���@tj�M�f���E�   �M��tX�}� t&�U�R�E�P�M����P�M�Q�U�R������E���E�P�M�Q�M��h���E��U��UЋE�P�M����E�V�T�}� t&�M�Q�U�R�M��@��P�E�P�M�Q�\�����E���U�R�E�P�M�����E��M��M��U�R�M�A���E^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���� ����u3���   ��   � ����0|8� ����9*� ����/�M�� ���� ��E��   �   �E�    � ����@tY� ����u3��k�7� ����A|$� ����P�U���� ���T
��U������2� ���� �뚋 ��� ���� ���@t�����E���]����������������������������������������������������������������������̋�U����   � ����?u� ��B��$tj�M����E�  � ���� ����U����E̋��M���\�������M���
���M���
����\������E����MЉ��M�������M�������E� � ����?u/� ���� ��U�Rj��T���P�y����P�M�������jj��L���Q�A�����P�M������M�������t�8��U���up��D���P������Pj<��<���Q������P�M������M��?���Ѓ�>u
j �M�����j>�M��y����E��t� ����t� ���� ��M����Ủ��E����M�Q�M�����E��]�����������������������������������������������������������������������������������������������������������������̋�U���|���3ŉE��E�   �M��*����9��M��i������  � �����  � ����@��  �}� t	�E�    �
j,�M��F���� ����0�U�x4�}�	.� ���� ��M�Q�U�R�������P�M��}����  � ��E�M������ ����Xu� ���� �htb�M������%  � ����$u7� ��H��$t)� ���� ��E�P��	����P�M��\�����   � ����?��   �E�P������������tkj�M�Q�M��)���U�R�����P�4����Eă}� t�E�P�M������.h�a�M�Q�U�Rh\b�E�P�L�����������P�M�������.h�a�M�Q�U�Rh\b�E�P���������d���P�M�������M��G���P�M�Q�L�����P�M��w���� �+U��~���e�����u�E�P��������M�Q�M������������9� �U�R�M�����E�M�3��U�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���  ���3ŉE� ���M�� ���� ��E�������������R��  �����������$�p��EP��������E�  � ����@u$� ���� �h|b�M�����E�S  �3��D���Q�A�����P�URh$_��L����X������.����E�  �EP�������E�
  �M�Q�N������U�R�B������M����������   �M�������t{jd�E�P�M��P�����uj�M�+����E�  �M��M��U���-u�E��E��E�.��E�.�M�Q�URje��4���P�M�Q��<����������R������m����E�]  �j�M������E�I  ��x���R������������tSj��h���P��x���������h���Q�����P�4�����d�����d��� t��d���R�M�����E��  �E���Du5h�a�MQ��x���Rh\b��,���P��������������E�  �3h�a�MQ��x���Rh8b��$���P�r������������E�m  �h  j j ��\���Q�T����������R��������\���P�M�<����E�/  j{��T����i����M�������������H|3������J~�(�����R�������P��T����
���j,��T��������E���������������F������������wx�������$��������P�������P��T�������j,��T����/��������Q�������P��T�������j,��T�������������R������P��T����c���j}�EP��T��������E�-�+� ���� �j�M�����E�j�M�t����E�M�3�������]Ë�5�����V��B�1���S� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �M��h���� ���E��M�����E��}���  uj�M�x����E�  �B�}���  u�EPj�MQ�'������E�  ��}���  u�UR�M������E�j  �E�% �  �0  �M��� �  t�U���   3���   ���������M��� `  ��Ƀ����������� t�U���   �� �����E�%   �� ����� ��� t>�M��� �  t�U���   3���   ���������
ǅ����    ������ ��
  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ t|�M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� �  t�U���   3���   ���������
ǅ����    ������ ��	  �M��� @  tM������t/�E�����t&�U�R�\�����Pj �E�P�i�����P�M��W�����M�Q�6�����P�M�������U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t�E�%   ��������M���   ������������ �-  �U��� �  t�E�%   3�=   ���������
ǅ����    ������ ��   �U�R�K�����P��|���Pj{�M�Q�M������������P�M������U�R�r������������u1h�c��l���P�M�Qj,��t���R�5������������P�M�����h�c�M��G����E�P�������������tR������tI������u@�M�Q��T���Rj ��\���P�M�Qj ��d���R����������������8���P�M������  �M��U����M��M����M��E����M��=����M��5����E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ �"  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t[�M���   ��   uJ��L���R�������P�M�������D���P�������P�M�������<���Q������P�M��m����k�U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� t'�E�%   =   u��4���Q�Q�����P�M�� �����,���R�9�����P�M�������E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t8�U��� �  t�E�%   3�=   ���������
ǅ����   ������ u;������t��$���R������P�M�����������P������P�M��w����e�����tO������t,�M�Q�����R�����P���������;���P�M�����������Q�m�����P�M��!����������R�S�����P�M������M�K�����uA�M��?�����u)� �����u �EPj ������Q�J�����P�M��������UR�M��*����E�    �M�������}� tNj ������P�/�����Ph�c������Q�d�����P�M�����������t�U�R�M�U����E��  �bj h �j������������������� t�������V����������
ǅ����    �������E��M�Q������R������P�M��e����E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t�M���   ��������U���   ������������ ��  �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� ��   �M���   ��   uzj,������R�E�P������Qj,������R�E�P������Qj,������R�E�Ph�c������Q��������������������������������������P�M�������   �U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� tB�E�%   =   u3j,������Q�U�Rh�c������P�"�����������P�M��<����h�c�M������h�c������Q�M��>���P�M�����j)��x���R������P�W�����Pj(������Q�P�����������P�M�������U��� �  t�E�%   3�=   ����������U��� `  ��҃������������� ��   �E�% �  t�M���   3ҁ�   ��������E�% `  ����������������� t:�M��� �  t�U���   3���   ���������
ǅ����   ������ u�M�Q�M�����������t��p���R������P�M���������h���P�j�����P�M������(�����t�}� t�M�Q�M������U�R�M������  �EP�M������M��� �  u.�U��� |  �� h  u�E�P�MQ��������E��	  �1  �U��� �  u,�E�% |  = p  u�M�Q�UR�~������E�	  ��  �E�% �  u]�M��� |  �� `  uLh�c�UR��X���P������P��P���Qj{��`���R�M�������������������E�N	  �  �E�% �  u.�M��� |  �� |  u�U�R�EP��������E�	  �[  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ thXc�M��f����  �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tL�M��� �  t�U���   3���   ���������
ǅ����    ������ thc�M�������   �M��� �  t�U���   3���   ����������M��� `  ��Ƀ������������� t�U���   ��������E�%   ������������ tI�M��� �  t�U���   3���   ���������
ǅ����    ������ th�b�M�������0�M��� �  u%�U��� |  �� x  u�E�P�M�����E�  �M��� �  t�U���   3���   ����|�����M��� `  ��Ƀ���|�����|��� t�U���   ��x�����E�%   ��x�����x��� ��   �M��� �  t�U���   3���   ����t����
ǅt���    ��t��� u:�M��� �  t�U���   3���   ����p����
ǅp���    ��p��� t#�M�Qh�c��H���R�������P�M�������E�P��@���Q�������P�M��c����U��� �  t�E�%   3�=   ����l�����U��� `  ��҃���l�����l��� �x  �������R  �E�% �  t�M���   3ҁ�   ��h�����E�% `  �������h�����h��� t[�M��� �  t�U���   3���   ����d����
ǅd���   ��d��� t!�M�Qh�b��8���R�������P�M��o����E�% �  t�M���   ��   �s  �U��� �  t�E�%   3�=   ����`�����U��� `  ��҃���`�����`��� t�E�%   ��\�����M���   ��\�����\��� �$  �U��� �  t�E�%   3�=   ����X�����U��� `  ��҃���X�����X��� t�E�%   =   ��   �M��� �  t�U���   3���   ����T�����M��� `  ��Ƀ���T�����T��� t�U���   ��   tU�E�% �  t�M���   3ҁ�   ��P�����E�% `  �������P�����P��� t2�M���   ��   u!�U�Rh�b��0���P�:�����P�M������������  �M��� �  t�U���   3���   ����L�����M��� `  ��Ƀ���L�����L��� tl�U��� �  t�E�%�   3Ƀ�@����H�����U���   3���   ����H�����H��� t&�M�Qh�b��(���R������P�M������Z  �E�% �  t�M���   3ҁ�   ��D�����E�% `  �������D�����D��� tp�M��� �  t�U����   3����   ����@�����M���   3ҁ�   ��@�����@��� t&�E�Ph�b�� ���Q�������P�M��N����   �U��� �  t�E�%   3�=   ����<�����U��� `  ��҃���<�����<��� tb�E�% �  t�M����   ��Ƀ���8�����U���   ��҃���8�����8��� t!�E�Ph�b�����Q�!�����P�M������U��� �  t�E�%   3�=   ����4�����U��� `  ��҃���4�����4��� t�E�%   ��0�����M���   ��0�����0��� t*�������u!�U�Rh�b�����P������P�M������M���   t!�U�Rh�b�����P�_�����P�M�������M�Q�M�Y����E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���x�E�    � ����_u�U��� @  �U�� ���� �� ����A�  � ����Z�  � ����A�E�� ���� ��U��� �  �U��E���t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M�U����U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U��E��E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E܋M܉M��;�U��� �  t�E�%?����E���M��������M؋U؉U���E���  �E��k  �E����Eԃ}���   �M��$��	�U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M̋ỦUЋEЉE����E���  �E��  �  � ����$��  �E� � ���� �� ���Uȃ}�R�]  �E����	�$��	�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  � ��Q��Pu� ���� �� ���� �� ���Eă}�Q��   �M���T	�$�@	� ���� ��:����  � ���� �� ����0|C� ����95� ��� ��D
ѣ �������E��M���   �M��E��-  ��E���  �7� ���� ������	  �E���  �E���  �E���  �E���  ��  �E���  � ���� ���  �E�� ���� �� ����0|� ����5~$� ����t	�E���  ��E���  �E��z  � ����0�E��M��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��M���t�U���    �U���E�%�����E��M����M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  � ���� ���  � ����0��  � ����8��  � ���U� ���� ��M�������M��U�U��E���0�E��}��?  �M��$��	�U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C� ����9u� ���� ��E���  �� ����t	�E���  ��E���  �E���]ÍI ����|���j���S�����'�>�U���j������� 																																																																					��������� �� 	� 	J	�	�	�		'	9	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j �������P�M������ ����tl� ���E� ���� ��U�U�}�0t�}�2t�}�5t(�5htb�M��P����&�E�P������P�M������j�M������E�(�
j�M��1���h�c�M������M�Q�M�O����E��]���������������������������������������������������̋�U���@�M��;���j j�E�P�������P�M��h����M��h�����uN� ����tA� ����@t4�U�R�E�Ph�a�M�Q�U�R�g��������������螾��P�M������ ����@u� ���� ��b� ����tj�M������J�M�������tj�M������2�U�R�E�Ph�a�M�Qj�M��������b���������P�M�莸���U�R�M�����E��]��������������������������������������������������������������������������̋�U���� �����  � ����A�E�� ���� ��}���   j�M�������e�������   �U�����U��}���   �E���
	�$��		j� �����P�M������|j�������P�M������gj�������P�M������Rj�������P�M��o����=j������P�M��Z����(j������P�M��E����j������P�M��0����U�R�M�����E� �j�M������E��j�M������E��]ÍI +		@		U		j				�		�		�		 ��������������������������������������������������������������������������������������������̋�U�� ����@u"� ���� ��EP�M�Y����E���MQ�UR�u������E]�����������������������̋�U��� �EP�M������ ���U��}� t�}�?tq�}�Xt��   �E�Pj�MQ�}������E��   � ���� ��M��v�����thtb�M�3����E�   ��E�Ph�c�MQ��������E�w� ���� ��E�k�j �M������P�E�P�M�Q�U�R迵����P�M��'����E�P�MQ�������E�$�U�R�M�����E��E�P�MQ轹�����E��]�������������������������������������������������������������������������̋�U���<�M��K���� ���Mȃ}�B��  �U���	�$� 	�MQj�UR�������E�j  h�c�M��O����M������u
j �M��V����EP�M������ ���� ��E�$_�U�R�M�����P�E�P�MQ��������E�   � ��B��$t<� ��Q��u�EPj�MQ�|������E��  �j�M�����E�  � ���� �� ���Mă}�T�o  �U���|	�$�X	� ���� ��UR�EP��������E�Y  � ���� �j�UR�EP�=������E�0  � ���� ��E�k�j �M�豼��P�U�R�EP�M�Q�q�����P�UR�������E��   ��   h�c�M�������M������u
j �M��Ͳ���EP�M������ ���� ��E��^�U�R�M�����P�E�P�MQ�n������E�z� ���� �j�M�8����E�\�G� ���� �h�c�M�Ѳ���E�;�&�MQj�UR��������E�"j�M������E��EP�MQ�������E��]Ë�v	�	�	�	�	 ��	z	�	�	<		�	�	�	 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� � ���M�}�XtD�}�Zt�`� ���� ��Դ����t	�E���E� d�E�P�M�w����E��   � ���� �htb�M�S����E��   �U�R�������M�蕶������   � ���M�}� t�}�@t`�}�Zt�v�U�R�M������E�   � ���� ��(�����t	�E��c��E��c�M�Q�U�R�M�����P�M�����E�>� ���� ��M�Q�M�z����E� j�M������E���U�R�M�X����E��]��������������������������������������������������������������������������������������������̋�U���,�E�   �M������M��Z������  � ����@��   � ����Z��   �}� t	�E�    �
j,�M��6���� ������   � ����0�M�x3�}�	-� ���� ��E�P�M�Q��輱��P�M��[����k� ��U�M��c���P�E�P�h������ �+M��~��芰����u�U�R�������E�P�M������ �;M�u
j�M�葱���j�M�萰���������U�R�M贿���E��]����������������������������������������������������������������������������������������̋�U���(� ����tg� ����Zu'� ���� ��M��R���P�M�����E�^�0j)�UR�E�P�t�����Phd�M�Q����������°���E�,�*j)�URj�E�Phd�M��������������蔰���E��]�������������������������������������������������������̋�U���x� �����k  � ���E�� ���� ��E� �E������M��f����U��U��E���C�E��}��   �M����	�$��	h�d�M������?  h�d�M��m����-  h�d�M��[����  h�d�M��I����	  h�d�M��7�����  h�d�M��%���h�d�M��E�����  �E����E���  � ���U��E�E�� ���� ��U��U��}�Y�8  �E���	�$��	�E������(  h�d�M�詸���  h�d�M�藸���  h�d�M�腸����   h�d�M��s�����   h�d�M��a�����   htd�M��O����   hhd�M��=����   h\d�M��+����   � ���� ��E�P�D�����P�M�������M��˹����t�M�Q�M�c����E�~  �R�UR�E�P�r�����PhTd�MQ�(������E�R  � ���� �j�M��ԭ���hHd�M�获���Qhtb�M������B� ���� ��M�Q蝳����P�M��P����M��$�����t�U�R�M輻���E��  �}����   �E��E��M���C�M��}���   �U���x	�$�h	�M�Qh<d�U�R�[�����P�M��ݨ���e�E�Ph0d�M�Q�;�����P�M�轨���E�U�U��E���E�E��}�w/�M����	�$��	�E�Ph<d�M�Q�������P�M��v����M�J�����u�URj �E�P�a�����P�M������M�Q�M�Ǻ���E��   ��   �M������UR�M�覺���}��uF�M������E�P�M�Q�U�R脸�����M��i�����uhL_�M������E�P�M�_����E�}�M誷����tA�M���t$h(d�M�������U���thd�M��ؿ����E���th�c�M�蔵���M�Q�U�R�EP詷�����E���MQj�UR� ������E��]�`	r	�	�	�	�	�	�	`	�	o	   










	�I 6		H	Z	l	~	�	6	*	�	�	�	Q	 	
��	�	&	k	 �I M	k	     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�������t�Q�����u	�E�   ��E�    �EЉE��M��C���� ���U̡ ���� ��M̉Mȃ}�Y��   �U����	�$�t	� ���� �h)e�M�ݤ���E�   h e�M��)����khe�M������\he�M������Mh e�M�������>h�d�M������/�����E��U�R�a�����Ph�d�E�P�/�����P�M�豣���M��c����}� t�M�Q�M�藣���U�R萦����P�M��!����E�P�M������E��]Ë��	�	�	�		�	�	0	 ���������������������������������������������������������������������������������������������������������������������������������̋�U��EP�u������E]����������̋�U����M������� ������   � ���E�M��0�M�}�wH�U��$��	hLe�M��
����>hDe�M�������/�-h<e�M������h�d�M��ۯ���j�M贶���E�~� ���M� ���� ��E�E�M��1�M�}�w/�U����	�$��	�M�Qh<d�U�R�߶����P�M��a����E�P�M�ٳ���E��j�M�4����E��]��	�	�	�	�	�			b	�	    ��������������������������������������������������������������������������������������������̋�U����   � ����u�URj�EP�L������E�  � ����6|� ����9~ � ����_tj�M�=����E��  � ����6�U�� ���� ��}�)u[� ����t2� ����=�M�� ���� ��}�|�}�~�E�������EPj�MQ薱�����E�M  ��}� |�}�~�E������}��uj�M蕴���E�   �M��O����UR�M������E����  �M�Qh�a�U�R�ݴ����P�M��_���� ����t5�U�R�E�P�M�Q聡����Pj �U�R�9�������谤��P�M�� �����E�Pj�M�Q�а����P�M������ ����t1� ����@u� ���� ��j�M迳���E�J  ��M�Qj�UR�w������E�.  �C�����t�E�P�,�����P�M�荞����M�Q������P�M������U���tS������t5�E�P�M�Q�U�R�>�����Pj �E�P�K��������£��P�M��2�����M�Q������P�M�諸��虢����t)�U�R��x���P�M�Q�Π�������{���P�M��������p���R譠����P�M��a����M襭����u.j)��`���P�M�Qj(��h���R谫����������P�M�藝��j h �j���������\�����\��� t��\����&�����0����
ǅ0���    ��0����E��M�Q�U�R�l�����j)��D���P��T���Q�'�����Pj(��L���R� ��������u���P�M�覣��蟥����t�E���t�M�Q�M�艣���?�����t��<���R�	�����P�M��h������4���P������P�M��?����}� t�M�Q�M�蝜���j�M聱���E��U�R�M�����E��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���� ������   � ����6|� ����9~� ����_un�UR�M�辛���M������u$�M�ܪ����u�M襭����u�EP�M�胡���M踪����u�MQ�M��k����U�R�EP�M������E�   �>j �MQ�UR�EP�M�Q�'������U�3Ƀ�*��Q�U�R�EP藝�����E�m�kj�M��X����MQ�M�蔲���M�0�����u�UR�M������M������u"�M������u
j �M��J����EP�M�赠���M�Q�M莬���E��]��������������������������������������������������������������������������������������������������̋�U���4�M��K���� ���� �� ���UЀ}�At�}�BtN�}�C��   �   �} u%�E����&u	�E�_��E��^�E�M̉� ���� ��  �} tj�M������E�}  �E� j>�M��u���� ���� ��N  �U�_� ���� ��3  � ����t� ��H��uj�M蔭���E�  �} tj�M�|����E��   � ����0��� ��Q�DЉE� ���� ��}�v/j,�M��ð���U�3�PR�M��~���P�M�Q�M�谝��P�M�� ���j>�U�R�M��w���P�M��	���� ����$u� ���� ��j^�E�P�M��B���P�M��ԗ��� ����t� ���� ��
j�M�������M�肶���M�Q�M�����E��M�G����E��]�����������������������������������������������������������������������������������������������������������������������������������������������������̋�U���$  �M�蘠���E� � �����  � ����$u8�MQ�U�R�EP�M�Q�������M��x�����u�U�R�M�����E�  � ��� ��3҃�A����+��+ʉM�M������M������E�   �E艅����������t������tw��������   �  藚����tW�c�����tN�M��ۥ����u/j�E�����P�M�Qj �U�R�M��C�����蛤��P�M��Ε���j������P�M��ģ���   �2�����tN�M�������u/j
������P�E�Pj �M�Q�M��������?���P�M��r����j
躞����P�M��h����`�ٙ����tN�M��&�����u/j	萞����P�U�Rj �E�P�M�莙��������P�M������j	�a�����P�M�������E�    �}� t|� ���� �� ����$u8�MQ�U�R�EP�M�Q�!������M�蔤����u�U�R�M�,����E�  � ��� ��3҃�A����+��+ʉM�}� �)���� ����t� ���� ��}���  �EP�M������M�Q�U�R�M�赙��P�M��%����M��������u)�E�P��|���Qj �U�R�M��e�����耙��P�M������M��ģ����u,�E�P��l���Qj ��t���R�M��-������H���P�M�踓���E���  �} tj�M茨���E�  �M���tz�E�Ph�a��d���Q������P�M��i���� ����t,�M�Q��T���R��\���P脕���������P�M��2�����M�Qj��L���R�ߤ����P�M������$� ����t��D���R�7�����P�M��|���� ����uj�M��#����/� ��� ���� ���@tj�M蝧���E�  �#�����t[�U��������������t�B�} tj�M�e����E�t  �E�P��4���Q��<���R�@��������ӗ��P�M��C����#�E����u��,���Q������P�M�讬���U��t!�E�Ph\e��$���Q�s�����P�M�������U��t!�E�PhTe�����Q�J�����P�M��̑���} ��   �M薡������   �M�[�����u�M�z�����t:�M������t�UR�M�肑����EPj �����Q�t�����P�M������@�UR������Pj �����Q�URj �����P�@�������蕕����谖��P�M�迗���*�M������u�MQj ������R������P�M�蓗���M�������E���t�M������M�Q�M�T����E��   �j�M謥���E�   �   �} ux�M�}�����ul�M�F�����u�M�e�����t�URj�EP�7������E�u�9�MQ�URj ������P�MQj������R�
�������褔����迕���E�:�8�} u%�M�������u�EPj�MQ�ѡ�����E��j�M�����E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���� �����  �} t]� ����XuO� ���� ��M�ʝ����thtb�M臎���E��   ��URh�c�EP�3������E��   � ����Yu%� ���� ��MQ�UR豗�����E�   �EP�M�Q� ������M�ǐ����t �U�Rhxe�E�P�Ǣ����P�M��I����*�M�r�����t�M�Qhhe�U�R蛢����P�M������E�P�M蕟���E���MQj�UR輞�����E��]��������������������������������������������������������������������������������̋�U���   � �����s  �ə���E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M�������������謐��P�MQ�������E�  �  �M��ߕ���M莝����thL_�M��D����M��Y�����tR�U��E����E���tB� ����t5j]�E�Pj �M�Q�-�����Pj[�U�R�ə����������P�M��O���뢋M肛����u^�M������t�E�P�M�Q�M����P�M��}����7�U�R�E�Pj)�M�Q�URj(�E�P�d�������蹏�����Ԑ��P�M��D����M�Q�U�R� ������M������E�P�M褝���E�   �   �M������uSj]��|���Qj�U�Rh�e�E�P�MQj(�U�R��������蚙����肪�����-���P�EP�h������E�?�=j]��d���Qj��l���Rj[��t����[������A���������P�EP�'������E��]��������������������������������������������������������������������������������������������������������������������������������������������������̋�U���j'�EPj �M�Q�#�����Pj`�U�R迗�����������E��]�����������������������̋�U����E�k�j�M��2���P�E�P�M��%���P�MQ�������E��]����������������������̋�U��Q�E�8_�E�P�MQ�UR�EP�g������E��]��������������������̋�U��Q�E�k��E�P�MQ�UR�EP�'������E��]��������������������̋�U��EP�MQ�UR�EP�������E]��������������̋�U��j�EP�ܛ�����E]��������̋�U��j �EP輛�����E]��������̋�U��j �EP蜛�����E]��������̋�U��EP�MQ�2������E]������̋�U��Q� ���M��}� t)�}�At�0� ���� �h�e�M聈���E�j�M踜���E�j�M詜���E��]���������������������������������̋�U���@�EP�M������M��ʖ�����b  � �����Q  �E�P�M�Qj �U�R�E�P�8�������蠋����軌��P�M��+����M��x������  � ����@��   h�e�M��4����M��I�������   � ������   � ����@txj'�M�Q�U�R�������Pj`�E�P趔����������P�M��<���� ����@u� ���� ��M��ϕ����t� ����@th�e�M�蓞���Z����M�裕����t � ����u
j�M�聉��j}�M��R���� ����@u� ���� ��'�M��X�����t�U�Rj�E�P豗����P�M������M�Q�M�\����E��]����������������������������������������������������������������������������������������������������������������̋�U��EP�4������E]����������̋�U����E�k�j �M�����P�E�P�M��Վ��P�MQ蝅�����E��]����������������������̋�U����EP�M��a���h�e�M������M�Q������P�M��Z���j}�M��ل��� ����@u� ���� ��U�R�M�����E��]��������������������������������̋�U���,j h �j胗�����E��}� t�M������E���E�    �EԉE�M�Q�U�R�m������EP�M�Qj �U�R�E�P���������Y������t���P�M������M�Q�M�\����E��]������������������������������������������������̋�U��0��������]����������̋�U��0�%   �����]��������̋�U��0��������]����������̋�U��0��������]����������̋�U��0��������]����������̋�U��0���`3Ƀ�`����]�������̋�U��0�%�   �����]��������̋�U��0�%   �����]��������̋�U��0�%   �����]��������̋�U��0�%   ]���������������̋�U��0�%    ]���������������̋�U��0�% @  ]���������������̋�U��0�% �  �����]��������̋�U��0�%   �����]��������̋�U���%�����t�E��`���M��`��]���������������������̋�U��0��������]����������̋�U��EP�MQ� �����]�������̋�U����M�E������E�} t�MQ�U��Ѓ���   ��   �} w�E   �M�Q;U��   �}   v3��   jh �h  �'������E��}� t�M��p����E���E�    �E��E��}� tA�M�y t�U�B�M���U�E��B��M�U��Q�E�M��H�   +U�E�P�3��!��M�Q+U�E�P�M�Q�E�H�D
��]� ���������������������������������������������������������������������̋�U��Q�M��E��     �E���]�������̋�U����EP�MQ�UR�M�蚖�����T����E��]���������������������̋�U����EP�MQ�UR�M�腔���������E��]����������������������̋�U����EP�MQ�UR�M��������Մ���E��]����������������������̋�U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]�����������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��i����E���]� ������������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��} tdj h �j�������E��}� t�EP�M��J����E���E�    �M��U��E����Ƀ�������   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ���������������������������������������������������������������������������������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t%�MQ��"  ���E��}� v�U�R�EP�M�蒍���E���]� ���������������������������������������������������������������������̋�U���V�M�E�H�� ����U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E�H�������U�J�E��     �M�Q�������E�P�M�Q�������E�P�M�Q�������E�P�M�Q������E�P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	�w����t�U����U���E�H�� ������U�J�   ������E�P�M�Q�M��,����U����t<�U�E���M�	���u�;�t�U�B% ������M�A�U��    �!�M���~����u�E�H�� ������U�J��E�H�� ������U�J��E�H�� ������U�J�E�^��]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��0�%   ]���������������̋�U���$���3ŉE��M܍E��E��M܋Q�� ����E܉P�M��    �U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%�����M܉A�U܋B%����M܉A�U�� �E����E�j j
�MQ�UR������0�� �M��j j
�UR�EP臒���E�U�MMu��U��E�+й   +�Q�U�R�M�菈���E܋M�3���v����]� ����������������������������������������������������������������������������������������̋�U���(���3ŉE��M؍E��E܋M؋Q�� ����E؉P�M��    �U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%�����M؉A�U؋B%����M؉A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U܃��U�j j
�EP�MQ�R�����0�� �U܈j j
�EP�MQ�ΐ���E�U�UUu��E��t�M܃��M܋U��-�E܍M�+��   +�R�E�P�M�迆���E؋M�3���t����]� ��������������������������������������������������������������������������������������������������������̋�U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP�F������M���U��: u�E��H�� ������U��J�E���]� �����������������������������������������������������������������������̋�U��Q�M��E��H����3�������]���������������̋�U��Q�M��E�3Ƀ8 ������]������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J�E���]��������������̋�U��Q�M��E��@������]�������̋�U����M��M��������u�E��H��	��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��M�謀����u�E��H��   �U��J��]���������������������̋�U����M��M��j�����u�E��H��
��t	�E�   ��E�    �E���]��������������������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��   �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H��    �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� @  �U��J��]�����������������̋�U��Q�M��E��@������]�������̋�U��Q�M��E��H�� �  �U��J��]�����������������̋�U��Q�M��M��~����t3���E���U����ȋ�Ћ�]�����������������̋�U��Q�M��M��L~����t2���E���U����ȋB�Ћ�]����������������̋�U����M�M��
~����uX�} u*�M��������Ej h ��EP�>������E��M��M�} t �U�E�L�Q�UR�M������E��E��  ��} t�M� �E��]� �������������������������������������������̋�U��Q�M��M��\}����t�E��EP�MQ�U���M��	��B�Ћ�]� ����������������������̋�U����M�E�P�M�����MQ�M��Em���U�R�M����E��]� ����������������������̋�U����M�E�P�M��^���MQ�M������U�R�M�F���E��]� �����������������������̋�U����M�E�P�M�����MQ�M��s���U�R�M��~���E��]� �����������������������̋�U����M�E�P�M��~���MQ�M��/����U�R�M�~���E��]� �����������������������̋�U����M�E�P�M��n~���MQ�M��+o���U�R�M�V~���E��]� �����������������������̋�U����M��} t_j h �j��~�����E��}� t�EP�M��R�M���|���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ������������������������������������̋�U����M��M��Cz����tb�E��tZ�M��z����t�MQ�M��G����?j h �j��}�����E��}� t�UR�M��K����E���E�    �E�P�M������E���]� ���������������������������������������������̋�U����M��M��y����tu�} to�E���te�M���y����t�UR�M��x���Kj h �j�:}�����E��}� t�EP�  ��P�MQ�M��Qx���E���E�    �U�R�M��Y����E���]� ������������������������������������������̋�U��Q�M��M���x����tG�M�Py����t�M�pp��P�M��l���(�M��1y����t�EP�M��Ei����M�R�M������E���]� ��������������������������̋�U����M��M��Sx������   �} ��   �M���x����t�EP�M��Mr���j�M��o����t�M��o����u@j h �j��{�����E��}� t�MQ�M��p���E���E�    �U�R�M������M�yo��P�M��k���E���]� ���������������������������������������������̋�U��Q�M��M��uw����tC�M���w����u�}t�}u�EP�M��:l����} u��MQ�ă����P�M��m~���E���]� ������������������������������̋�U����M��M��n����t3�M��v����u'�M�n���E��E�%�   �M��Q�� ���ЋE��P�E���]� ���������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��iy���E���]� ������������������������������������������������������������̋�U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�  ��P�UR�M��Vx���E���]� ���������������������������������������������������������̋�U��Q�M��E��M���I�H�E���]� �������������̋�U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj h �j�_w�����E��}� t�MQ�M��k���E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������̋�U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ�~�����U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ������������������������������������������������������������������̋�U����M�E�8 tj�M��Vf���  �} ��   �} ��   �M�M��}� t�}�t�u�U�B% ������M�A�   j h �j��t�����E��}� t�U�P�M��Pz���E���E�    �M�U��E�8 u�M�Q�� ������E�P�[j h �j�t�����E��}� t�MQ�UR�M��o���E���E�    �E�M��U�: u�E�H�� ������U�J��E�H�� ������U�J��]� ����������������������������������������������������������������������������������������̋�U��Q�M��E�3Ƀ8	������]������̋�U��Q�M��E�� �����E���]�������̋�U����M�M��Uc����uf�M�p����uZj h �j�hs�����E��}� t�EP�M��r���E���E�    �M��M��}� t�U����M��U��M�U��T��E��]� �����������������������������������������̋�U��Q�M��} |�}	~j�M�t���E�;�9�E��8�t
�M��U;~j�M�_t���E���E�M��T�R�M��q���E��]� ��������������������������̋�U��Q�M��E�� �e�E���]�������̋�U��Q�M��M��x���E�� �e�M��U�Q�E���]� �������������������̋�U��Q�M��   ��]��������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E;Es�M�U��B��M���M�E��]� �����������������̋�U����M��M���w���E�� �e�} tP�} tJj h ��MQ�Qq�����E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ�S  ����U��B    �E��@    �E���]� ������������������������������������������������̋�U��Q�M��E��@��]�������������̋�U����M��E��x t�M��Q�E��H�T
��U���E� �E���]����������������������������̋�U��Q�M��E��HQ�U��BP�MQ�UR�{������]� ������������������̋�U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�"  ���EE��]���������������������̋�U����M��M��7v���E�� �e�} t#�M�oc����t�M�bc����u	�E�    ��M�M��U��E��B�E���]� ����������������������������������̋�U����M��E��x t�M��I��x���E���E�    �E���]��������������̋�U����M��E��x t�M��I�u���E���E� �E���]�����������������̋�U����M��E��x t�MQ�UR�E��H�s���E���M�M��E���]� ��������������������̋�U��Q�M��M���t���E�� �e�M��U�Q�E��H����Ƀ�����U��J�E���]� ��������������������������̋�U��Q�M��E��@��]�������������̋�U��Q�M��E��x��,"�e��]�����������������̋�U��Q�M��E��xujh�e�MQ�UR�y������E��]� ���������������������������̋�U��j�h�.d�    P���3�P�E�d�    �����uM���������E�    j ����_��j����_��j�����^��j�����^���E������} |�}}�Ek��������M�d�    Y��]��������������������������������������������������������̋�U��Q�M��M��	s���E�� �e�M��U�Q�E��M�H�U��B�����E���]� ����������������̋�U��QV�M��E��x }.�M��Q�E��H���Ћ��M��Q�E��H������M��q�U��B^��]��������������������̋�U����M��E��H�U��B��ȋB�ЈE��M���u�U��B�M��I��B�ЈE��E���]������������������������̋�U����M��EP�MQ�U��B�M��I��B�ЉE��M�;Ms�UR�E�P�M��Q�E��H��B�����E���]� ����������������������̋�U��Q�E�    �	�E���E�M���t�E����E���E���]����������������������������̋�U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]��������������������������̋�U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]������������������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uh�fj jEh8fj�]������u̃}� u.�et���    j jEh8fhfh�f�pn��������  �MQ�M��f���} �  �M��\����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M��ot���E��O  �M����M��U���U뱋E��EԍM��Et���E��%  �  �MQ�URj��EPj	�M��[����QR��E��}� t�E����EЍM���s���E���  ����zt*�Vs��� *   3ɋUf�
�E������M���s���E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M���Z��P�M��R��\������t@�E��H��u,��r��� *   3ҋEf��E������M��Cs���E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M��{Z����QR��E��}� u*�br��� *   3��Mf��E������M���r���E��   �U��U��M��r���E��   �   �M��Z��� �x u�MQ�]�����E��M��r���E��j�`j j j��URj	�M���Y��� �HQ��E��}� u!��q��� *   �E������M��=r���E�� ��U����U��M��%r���E���M��r����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�UR�EP��^����]�����������������̋�U��=�� uhH��EP�MQ�UR�$S������j �EP�MQ�UR�
S����]�����������������������������̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!hXgj h�   h8fj�FX������u̃}� u3�o���    j h�   h8fh4ghXg�i�����   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R�4X�����} t	�E�     �MQ�M��la���U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h gj h  h8fj�DW������u̃}� u@�n���    j h  h8fh4gh g�h�����E�   �M���n���E���  �M��aV��P�E�P�MQ�UR��\�����E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P� W������m����MЍM��`n���E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9��s����M��	�U���U��E���Ph�   �M��Q�dV�����U�9U����E�u!h�fj h  h8fj�U������u̃}� u=�m��� "   j h  h8fh4gh�f�g�����E�"   �M��gm���E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM��,m���Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�l����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�j jh�hj��S������u̃}� u0�-k���    j jh�hh�hh��8e�����   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�S����3҃} �U��}� uhL�j jh�hj�S������u̃}� u0�hj���    j jh�hh�hhL��sd�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���M܋U�Rh�   �E��P��R�����hh��t3�t	�E�   ��E�    �E؉E�}� uhhj j h�hj��Q������u̃}� u0�]i���    j j h�hh�hhh�hc�����   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���MԋU�Rh�   �E��P�Q��������t3�t	�E�   ��E�    �EЉE�}� uh��j j*h�hj��P������u̃}� u-�Oh��� "   j j*h�hh�hh���Zb�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9��s����U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR��P����3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uht�j jphP�j��N������u̃}� u.�Of���    j jphP�hDiht��Z`��������R  �} t�} u	�E�    ��E�   �M̉MЃ}� uh�j jshP�j�tN������u̃}� u.��e���    j jshP�hDih���_���������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �_�����Eă}��t�E���UU�B� �E��x }�����������]��������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh(��I�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh(��H�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h�ij h�   hP�j��K������u̃}� u1�Ic���    j h�   hP�h�ih�i�Q]���������  �} t�} v	�E�   ��E�    �U�U�}� u!hpij h�   hP�j�hK������u̃}� u1��b���    j h�   hP�h�ihpi��\��������d  �MQ�UR�EP�MQ�URh:��YG�����E��}� }U�E�  �}�tI�}���t@�}v:�M��9��s����U��	�E���E�M�Qh�   �U��R�8K�����}��uu3�t	�E�   ��E�    �M�M��}� u!hj h�   hP�j�kJ������u̃}� u.��a��� "   j h�   hP�h�ih��[��������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9��s
����E���M����U+щU��E�Ph�   �M��U�D
P�VJ�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�i]����]���������������̋�U���,�E������E�    3��} ���E�}� u!h�ij h  hP�j�H������u̃}� u1�`���    j h  hP�hjh�i�Z��������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!hpij h  hP�j�H������u̃}� u1�y_���    j h  hP�hjhpi�Y��������|  �M;M��   �<_����U��EP�MQ�UR�E��P�MQh:���C�����E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9��s����U���E���M+ȉM�U�Rh�   �E�M�TR��G�����^���8"u
�^���M������  �`�^����U��EP�MQ�UR�EP�MQh:��<C�����E��UU�B� �}��u"�}�u�A^���8"u
�7^���M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q��F�����}��uu3�t	�E�   ��E�    �E܉E�}� u!hj hB  hP�j�F������u̃}� u.�y]��� "   j hB  hP�hjh�W������������z�}�t\�}���tS�U���;UsH�E����M+�9��s����U���E����M+ȉM؋U�Rh�   �E��M�TR�F�����}� }	�E�������E��EԋEԋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�&=����]�����������̋�U����EPj �MQ�UR�EPh��l@�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh��
@�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uhl�j jfh@kj��B������u̃}� u0�CZ���    j jfh@kh0khl��NT�����   ��  3�;U��؉E�uhkj jgh@kj�B������u̃}� u0��Y���    j jgh@kh0khk��S�����   �  �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���UԋE�Ph�   �M��Q�{B����3҃} ��;U��؉E�uh�jj jih@kj�A������u̃}� u0� Y��� "   j jih@kh0kh�j�+S�����"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uhdjj jjh@kj�CA������u̃}� u0�X���    j jjh@kh0khdj�R�����   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!h0jj h�   h@kj�9@������u̃}� u0�W��� "   j h�   h@kh0kh0j�Q�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ������]�����������������̋�U��j �EP�MQ�UR�EP�T���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!hl�j h>  h@kj�=������u̃}� u3�U���    j h>  h@kh�khl��"O�����   �,  3�;U���؉E�u!hkj h?  h@kj�Q=������u̃}� u3�T���    j h?  h@kh�khk�N�����   ��  �U�� �}��tI�}����t@�}�v:�EЃ�9��s����M��	�UЃ��ŰE�Ph�   �Mԃ�Q�I=����3҃} ��;U���؉E�u!h�jj hA  h@kj�<������u̃}� u3��S��� "   j hA  h@kh�kh�j��M�����"   ��  �}r�}$w	�E�   ��E�    �UȉU܃}� u!hdjj hB  h@kj�<������u̃}� u3�iS���    j hB  h@kh�khdj�qM�����   �{  �E�    �MԉM��} t+�U��-�E����E��M����M��U�ڋE�� �؉U�E�M��M�U3�PR�MQ�UR�S���E�E3�QP�UR�EP�Q���E�U�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} w�} v�U�;U�r��E�;E�rl�M�� �U�;U���؉E�u!h0jj hf  h@kj��:������u̃}� u0�0R��� "   j hf  h@kh�kh0j�8L�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�B���]����������������̋�U���x���3ŉE��E�    �E�    �} t�} u3��  3��} ���EЃ}� uhplj jfh�kj��8������u̃}� u.�(P���    j jfh�kh�khpl�3J��������8  �UR�M��`B���} �.  �M���7��� �x ��   �M�;Msp�U�=�   ~"�O��� *   �E������M��2P���E���  �MM��U���M��E���E��u�M��M��M���O���E��  �U����U�눋E��E��M���O���E��  �  �M��97������   ��   �} v�UR�EP�  ���E�M�Qj �UR�EP�MQ�URj �M���6��� �HQ���E��}� t3�}� u-�UU��B���u	�M����M��U��U��M��>O���E���  �N��� *   �E������M��O���E���  ��  �E�Pj �MQ�URj��EPj �M��d6����QR���E��}� t�}� u�E����E��M���N���E��j  �}� u����zt"�N��� *   �E������M��N���E��7  �M�;M�  �U�Rj �M���5��� ���   Q�U�Rj�EPj �M���5����QR���E�}� t�}� t"�M��� *   �E������M��N���E���  �}� |�}�v"�yM��� *   �E������M���M���E��  �E�E�;Ev�M��M��M���M���E��t  �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M��zM���E��  벋U���U������E��E��M��TM���E���   ��   �M��4����y ur�E�    �U�U��	�Eȃ��EȋM����t;�E�����   ~"�vL��� *   �E������M���L���E��   �Ũ��U�벋ẺE��M���L���E��t�j�M�Qj j j j��URj �M��4��� �HQ���E��}� t�}� t��K��� *   �E������M��vL���E���U����U��M��`L���E���M��SL���M�3���.����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�������������������������������������̋�U��EP�MQ�UR�EP��E����]�����������������̋�U��j �EP�MQ�UR��E����]�������������������̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!h�lj h@  h�kj��1������u̃}� u3�'I���    j h@  h�kh�lh�l�/C�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�1�����} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h gj hL  h�kj��0������u̃}� u3�5H���    j hL  h�kh�lh g�=B�����   �  �MQ�U�R�EP�MQ�D�����E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U؋E�Ph�   �M��Q�0�����G��� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���MԋU�Rh�   �E��P�0�����M9M���ډU�u!h�lj hd  h�kj�f/������u̃}� u0��F��� "   j hd  h�kh�lh�l��@�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�MQ�C.����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�j jh�hj�-������u̃}� u0�E���    j jh�hh�mh��(?�����   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R�-����3��} ���E��}� uhL�j jh�hj��,������u̃}� u0�TD���    j jh�hh�mhL��_>�����   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E܋M���Qh�   �U��R�,�����hh��t3�t	�E�   ��E�    �U؉U�}� uhhj j h�hj��+������u̃}� u0�DC���    j j h�hh�mhh�O=�����   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���MԋU���Rh�   �E��P�+��������t3�t	�E�   ��E�    �EЉE�}� uh��j j*h�hj��*������u̃}� u-�0B��� "   j j*h�hh�mh���;<�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9��s����U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR�*����3���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!ht�j h�   h�mj��(������u̃}� u1�,@���    j h�   h�mh�mht��4:��������  �} t�} u	�E�    ��E�   �M̉MЃ}� u!h�j h�   h�mj�K(������u̃}� u1�?���    j h�   h�mh�mh��9��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �K9�����Eă}��tY�U��B���E��M��U��Q�}� |"�E��� 3ҁ��   �U��E�����U��
��E�Pj ��8�����E��}��t�E�� 3ɋU�Ef�LP��M��y }�����������]��������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EPj �MQ�UR�EPh���00�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQh����/�����E��}� }	�E�������U��U��E���]������������������������̋�U��� �E�����3��} ���E��}� u!h�ij h  h�mj�8%������u̃}� u1�<���    j h  h�mh�nh�i�6���������  �} t�} v	�E�   ��E�    �U�U�}� u!hPnj h  h�mj�$������u̃}� u1�<���    j h  h�mh�nhPn�!6��������j  �MQ�UR�EP�MQ�URh���}.�����E��}� }X3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M�U���Rh�   �E��P�$�����}��uu3�t	�E�   ��E�    �U�U��}� u!hj h  h�mj�#������u̃}� u.�;��� "   j h  h�mh�nh�!5��������m�}� |d�}�t^�}���tU�M���;MsJ�U����E+�9��s����M���U����E+E��M���Qh�   �U��E�LPQ�#�����E���]���������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�C*����]���������������̋�U���,�E������E�    3��} ���E�}� u!h�ij h9  h�mj�"������u̃}� u1�b9���    j h9  h�mh�nh�i�j3��������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!hPnj h?  h�mj�h!������u̃}� u1��8���    j h?  h�mh�nhPn��2��������  �M;M��   �8����U��EP�MQ�UR�E��P�MQh���+�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9��s����U���E���M+ȉM�U���Rh�   �E�M�TAR�!������7���8"u
��7���M�������  �c��7����U��EP�MQ�UR�EP�MQh���Z*�����E�3ҋE�Mf�TA��}��u"�}�u�7���8"u
�~7���U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�) �����}��ux3�t	�E�   ��E�    �U܉U�}� u!hj hf  h�mj�\������u̃}� u1�6��� "   j hf  h�mh�nh��0��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9��s����M���U����E+E؋M���Qh�   �U��E�LPQ�B�����}� }	�E�������U��UԋEԋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�EP�MQ�(����]�����������̋�U����EPj �MQ�UR�EPhF��p'�����E��}� }	�E�������M��M��E���]��������������������������̋�U����EP�MQ�UR�EP�MQhF��'�����E��}� }	�E�������U��U��E���]������������������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�@   �E��j �MQ�UR�EP�MQ�$   �E��E���]��������������������������̋�U���03��} ���E�}� uhl�j jfh@kj�������u̃}� u0�s3���    j jfh@kh�nhl��~-�����   �  3�;U��؉E�uhkj jgh@kj�������u̃}� u0�3���    j jgh@kh�nhk�-�����   �  3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���EԋM���Qh�   �U��R�����3��} ����;E��ىM�uh�jj jih@kj��������u̃}� u0�L2��� "   j jih@kh�nh�j�W,�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uhdjj jjh@kj�o������u̃}� u0��1���    j jjh@kh�nhdj��+�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!h0jj h�   h@kj�\������u̃}� u0�0��� "   j h�   h@kh�nh0j��*�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�e�����]�����������������̋�U��j �EP�MQ�UR�EP�4���]������������������̋�U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�   ��]�����������������������̋�U���8�UЉM�3��}� ���E�}� u!hl�j h>  h@kj��������u̃}� u3�*.���    j h>  h@kh ohl��2(�����   �A  3�;U���؉E�u!hkj h?  h@kj�a������u̃}� u3��-���    j h?  h@kh ohk��'�����   ��  3ҋE�f��}��tK�}����tB�}�v<�MЃ�9��s����U��	�EЃ��E̋M���Qh�   �Uԃ�R�U����3��} ����;E���ىM�u!h�jj hA  h@kj�������u̃}� u3��,��� "   j hA  h@kh oh�j��&�����"   �  �}r�}$w	�E�   ��E�    �EȉE܃}� u!hdjj hB  h@kj�������u̃}� u3�u,���    j hB  h@kh ohdj�}&�����   �  �E�    �UԉU��} t0�-   �M�f��U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ�,���E�U3�PR�MQ�UR�*���E�U�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} w�} v�M�;M�r��U�;U�rn3��M�f��U�;U���؉E�u!h0jj hf  h@kj��������u̃}� u0�3+��� "   j hf  h@kh oh0j�;%�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�U�M�"���]����������������̋�U����  ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M�����E�    �%)���E�3Ƀ} �������������� u!h�j h  h��j�}������u̃����� uF��(���    j h  h��hoh���"����ǅ<��������M��1)����<����  3��} �������������� u!ht�j h  h��j��������u̃����� uF�S(���    j h  h��hoht��["����ǅ8��������M��(����8����!  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U����  ������ ��  �������� |%��������x��������H�����,����
ǅ,���    ��,������������������������h�����������������(�����(����*  ��(����$��	�E�   ������Q�UR������P�h  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ��������$�����$����� ��$�����$���wL��$�����<�	�$�$�	�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�$�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP�#�����Ẽ}� }�E�������M�k�
�������DЉE��  �������� ����� �����I�� ����� ���.�  �� �����d�	�$�P�	�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  ���������	�$���	�M���0  u	�U��� �U��E�   �EP��!����f�������M��� tW���������   ������ƅ���� �M�����P�M������ ���   Q������R������P�<"������}�E�   �f������f�������������U��E�   �  �EP�V!���������������� t�������y u� ��U��E�P�������E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ����������������MQ� �����E��U��� ��   �}� u� ��E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M��d
��P�������Q�/������t������������������������������d�}� u	���M��E�   �U���|�������������������������t��|������t��|�������|����ɋ�|���+U����U��  �EP�������x����������   3�tǅ���   �
ǅ���    �������t�����t��� u!h�j h�  h��j��	������u̃�t��� uF�F!���    j h�  h��hoh��N����ǅ4��������M��!����4����  ��  �M��� t��x���f������f����x�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  h��j�Ḿ�]  Q������E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M�����P�U�R�E�P������Q�U�R�E�P��h���Q�H�R�l�Ѓ��E�%�   t%�}� u�M����P�M�Q�T�R�l�Ѓ���������gu)�M���   u�M��p��P�U�R�P�P�l�Ѓ��M����-u�E�   �E��M����M��U�R��
�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�h������X�����\����   �U���   t�EP�@������X�����\����   �M��� tB�U���@t�EP����������X�����\�����MQ�����������X�����\����=�U���@t�EP��������X�����\�����MQ�����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R������0��d����E��RP��T���P��P���Q�W����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �]  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M�����P�M���������   R��H���P������Q�9������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�  �������� |$�U���t������P�MQ��L���Rj �  ���}� tj�E�P�������E�    �"�����������0����M������0����M�3�������]Ð��	�	�	��	ָ	�	%�	`�	b�	m�	W�	L�	{�	��	 �I ��	D�	b�	O�	[�	 ��	��	�	�	M�	2�	��	��	#�	'�	ٿ	��	п	�	��	   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U���@�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!ht�j h�   h�mj�+�������u̃}� u1����    j h�   h�mh4oht����������V  3Ƀ} ���MЃ}� u!hj h�   h�mj���������u̃}� u1�"���    j h�   h�mh4oh�*���������   �E��@B   �M��U�Q�E��M��U��B����EP�MQ�UR�E�P������E��} u�E��   �M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj �������EȋE��H���MċU��EĉB�}� |!�M��� 3�%�   �E��M�����E����M�Qj ������E��E���]��������������������������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�I����]�������������������̋�U��EP�MQ�UR�EP�����]�����������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!ht�j h�  h�mj�[�������u̃}� u.����    j h�  h�mhToht���	��������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQh�������]������������������̋�U��EP�MQ�URh��������]����������������̋�U��EPj �MQhF������]������������������̋�U��EP�MQ�URhF��|����]����������������̋�U���@���3ŉE��E�    �w����E��E�    �E�    �E�    �=�� ��   h�� �Eԃ}� u3��  h�o�E�P�T�E��}� u3��  �M�Q�����h��U�R�TP�����h��E�P�TP�����h�o�M�Q�T�E��U�R������=�� tht�E�P�TP��������;M�th���;U�t]���P�l�EЋ��Q�l�Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W���;M�t���R�l�Eȃ}� t�UȉE�}� t*���;E�t ���Q�l�Eă}� t
�U�R�UĉE���P�l�E��}� t�MQ�UR�EP�M�Q�U���3��M�3��p�����]������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uht�j jphP�j���������u̃}� u.�?���    j jphP�h�oht��J��������   3Ƀ} ���MЃ}� uhj juhP�j�z�������u̃}� u.��
���    j juhP�h�oh����������   �E��@����M��AB   �U��E�B�M��U��EP�MQ�UR�E�P�������E��} u�E��Q�M��Q���ŰE��M̉H�}� |"�U���  3Ɂ��   �MȋU�����M����U�Rj ������EȋE���]������������������������������������������������������������������������������������������������������������̋�U��EPj �MQ�UR�
����]�������������������̋�U���,�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!ht�j h�  hP�j��������u̃}� u.�	���    j h�  hP�h�oht����������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]������������������������������������������������������̋�U��EPj �MQh(�������]������������������̋�U��EP�MQ�URh(�������]����������������̋�U��EPj �MQh��W�����]������������������̋�U��EP�MQ�URh��%�����]����������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    j�������E�    �EP�	����f�E��E������   �j�o������f�E�M�d�    Y_^[��]���������������������������������������������̋�U��Q�=���u�+����=���u���  �(j �E�Pj�MQ���R�H��u���  �f�E��]��������������������������������̋�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M������M��7�������   t1�M��$���� ���   thxpj jGh pj��������u̍M��������z u*�} t�Ef��Uf�
�E�   �M��V���E��R  �M�����P�E�Q����������   �M���������   ~R�M������ �M;��   |=3҃} ��R�EP�M��c�������   R�EPj	�M��L�����QR���uB�M��4���� �M;��   r�U�B��u"���� *   �E������M�����E��   �M����������   �U�M��l���E��k�a3��} ��P�MQj�URj	�M������ �HQ���u���� *   �E������M�����E���E�   �M��	���E���M�������]��������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�>����]�������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �}�u�0����     �	   �;  �} |�E;h�s	�E�   ��E�    �MԉM��}� uh�j j7h�qj��������u̃}� u;������     ���� 	   j j7h�qh�qh��������	   �  �E���M���������D
������؉E�uhj j8h�qj�*�������u̃}� u;�B����     ���� 	   j j8h�qh�qh�������	   �'  �} |�} r	�E�   ��E�    �UЉU؃}� uhtqj j9h�qj��������u̃}� u;�����     �����    j j9h�qh�qhtq�������   �   �MQ�������E�    �U���E���������T��t�EP�MQ�UR��������E��43�uh��j jAh�qj���������u��Y��� 	   �E�	   �E������   ��UR�#�����ËE�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���HV�E�    �E�    �E�    jj j �EP�������E؉U܋M�#M܃��t#jj j �UR�t������EЉUԋE�#Eԃ��u� ��� �  �M+MЋUUԉM�U�}� �?  
�}� �3  h   j��P�T�Eȃ}� u%�����    �E�   �E������E�������   h �  �EP�"������E�}� |	�}�   r	�E�   ��M�MċUĉU�}� |	�}�   r	�E�   ��E�E��M�Q�U�R�EP��������E�}��u(������8u�����    �E�   �E���E��U��*�E���M�+ȋE�M�E�}� �W���|
�}� �K����M�Q�UR�Z������E�Pj ��P�d�   �}� ~|�}� svj �MQ�UR�EP��������E��U��M�#M����tO�UR�������P������؃���E��U��E�#E����u!�C����    �E�   ����������0�M�#M����t'j �U�R�E�P�MQ�W������E��U��U�#U����u	������ �3�^��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�RP�EP�r������E��E������]����������̋�U��j�h8�h9�d�    P���SVW���1E�3�P�E�d�    �}�u�����     ����� 	   ����  �} |�E;h�s	�E�   ��E�    �M؉M��}� uh8�j jAh0rj���������u̃}� u9�����     �O���� 	   j jAh0rhrh8��Z���������/  �E���M���������D
������؉E�uh��j jBh0rj�s�������u̃}� u9�����     ������ 	   j jBh0rhrh�������������   �UR�v������E�    �E���M���������D
��t�MQ�UR�EP��������E��?�O���� 	   ������     �E�����3�uh��j jMh0rj��������u��E������   ��EP�������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP��������E��}��u5�4���� 	   3�uh�rj jjh0rj��������u̃���   �EPj �MQ�U�R���E��}��u���E���E�    �}� t�E�P�v���������;�M���U���������L����U���E���������L�E���]���������������������������������������������������������̋�U��j�hX�h9�d�    P���SVW���1E�3�P�E�d�    �} @  t-�} �  t$�}   t�}   t�}   t	�E�    ��E�   �EԉE��}� uhxsj j6h sj�A�������u̃}� u.�����    j j6h sh�rhxs����������  �}�u�n���� 	   ����  �} |�U;h�s	�E�   ��E�    �EЉE܃}� uh8�j j8h sj��������u̃}� u.�
���� 	   j j8h sh�rh8�����������  �U���E���������T������ډU�uh��j j9h sj�.�������u̃}� u.����� 	   j j9h sh�rh������������   �MQ�<������E�    �U���E���������T��t�EP�MQ�������E��4����� 	   3�uh��j jDh sj��������u��E������E������   ��MQ�������ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���M���������D
%�   �E��M���U���������L$�����щU��E�E�}�   $�}�   �a  �}� @  tm�}� �  t$�  �}�   �=  �}�   ��   �  �M���U���������L������U���E���������L�`  �E���M���������D
�   �M���U���������D�U���E���������T$�​E���M���������T$��   �M���U���������L�ɀ   �U���E���������L�E���M���������D
$$��M���U���������D$�u�U���E���������T�ʀ   �E���M���������T�M���U���������L$�က��U���E���������L$�}� u� �  ��}� u	� @  ���   ��]����������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} @  t�} �  t�}   t	�E�    ��E�   �E��E��}� u!h�tj h�   h sj�J�������u̃}� u0�����    j h�   h sh�th�t�������   ��URh ���3���]�����������������������������������������������������̋�U��Q3��} ���E��}� u!hXuj h�   h sj��������u̃}� u0������    j h�   h sh<uhXu��������   ��U� ��3���]���������������������������������̋�U���@�} �!  �EP�M������3Ƀ} ���M�}� uh �j j;h�uj���������u̃}� u=�=����    j j;h�uh�uh ��H������E�����M������E��  3��} ���E��}� uhL�j j<h�uj�i�������u̃}� u=������    j j<h�uh�uhL���������E�����M��&����E��1  ����;U����E�uh�uj j=h�uj���������u̃}� u=�W����    j j=h�uh�uh�u�b������E�����M������E��   �M�������z u)�EP�MQ�UR��������E̍M��|����E��   �m�E��MčM������P�U�R�m������E��E���E�M��U��M�����P�E�P�C������E��M���M�U���Ut�}� t�E�;E�t��M�+M��MȍM�������E��3���]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����=�� �Y  3��} ���E��}� u!h �j h�   h�uj��������u̃}� u3�s����    j h�   h�uh@vh ��{����������  3҃} �U��}� u!hL�j h�   h�uj��������u̃}� u3�����    j h�   h�uh@vhL������������   ����;M҃��U�u!h�uj h�   h�uj�:�������u̃}� u0�����    j h�   h�uh@vh�u�����������.�MQ�UR�EP�@�������j �MQ�UR�EP��������]��������������������������������������������������������������������������������������������������������̋�U��=�� uj �EP�MQ�URhH��:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�h�.d�    P��H���3�P�E�d�    �EP�M������E�    �} t�M�U�3��} ���Ẽ}� uhDwj j^h�vj��������u̃}� uD������    j j^h�vh�vhDw��������E�    �E������M��H����E��  �} t�}|�}$~	�E�    ��E�   �U��Uȃ}� uhXvj j_h�vj���������u̃}� uD�]����    j j_h�vh�vhXv�h������E�    �E������M������E��v  �M�M��E�    �U���E�M����M��M��������t0�M����������   ~�M������Pj�E�P�]������E��j�M�Q�M�����P�������E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} |�}t�}$~.�} t�U�E��E�    �E������M������E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M����M��U���E�M����M�����3��u�E�j�U�R�M��9���P��������t�E��0�E��Qh  �M�Q�M�����P�h�������t0�U��a|�E��z�M�� �M���U�U��E���7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M���U�E����E��!����M����M��U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4����� "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U���E��t�M��ىMЋUЉU��E������M��7����E��M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�������]���������������̋�U��=�� uj�EP�MQ�URhH���������j�EP�MQ�URj �n�����]�������������������������̋�U��j�EP�MQ�UR�EP�4�����]���������������̋�U����E�    �E�E�}� |,�}�~�}�t�����M��U����y����E��o3�t	�E�   ��E�    �U��U��}� uhxj j9h�wj��������u̃}� u+�����    j j9h�whdwhx�����������E���]���������������������������������������������������̋�U��E���]�����������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh�j jh�Fj��������u̃}� u0�����    j jh�FhHxh��������   �`  �} u`3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E�M���Qh�   �U��R������3���  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�;�����3Ƀ} ���M��}� uhL�j jh�Fj��������u̃}� u0������    j jh�FhHxhL���������   �2  �E�E��M�M��}�u7�U��Ef�f�
�U���M����M��U���U��t�E����E�t���}������t&�M;Mrh�j j+h�Fj���������u̋E��Mf�f��E���U����U��E���E��t�M����M�t�U���Ut���} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �E  3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E܋M���Qh�   �U��R����������t3�t	�E�   ��E�    �U؉U�}� uh��j j>h�Fj���������u̃}� u-�#���� "   j j>h�FhHxh���.������"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9��s����M���U+U����E+EԋM���Qh�   �U+U��E�LPQ������3���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�    �0���t
j
������������E��}� t
j�c������0���tjh  @j�������j�*�����]��������������������������������̋�U��Q�0��E��M��#M��U#Uʉ0��E���]���������������������̋�U����EP�M������MQ�UR�EP�MQ�M�����P�.   ���E�M������E��]�������������������������̋�U����E�    �E��Q�U�j j �EP�MQ���E�}� u3���   �}� ~63�u2�����3��u��r#h��  �E�L Q������P�������E���E�    �U�U��}� u3��s�E�P�M�Q�UR�EP����u�H�F�} uj j j j j��M�Qj �U�R���E��!j j �EP�MQj��U�Rj �E�P���E��M�Q��������E���]��������������������������������������������������������������������������̋�U���$�} t�} v	�E�   ��E�    �E�E��}� uh�j jh�xj�L�������u̃}� u0�����    j jh�xh`xh��������   �(  �E�    �U�U�} tI�E���t?�U����U��E�;Er�  �M�Uf�f��M���M��:   �E�f��M���M�U�U��}� ��   �E������   �U����U��E�;Er��  �M�U�f�f��M���M�U����U��E����uU����U��E����/t5�U����\t*�M����M��U�;Ur�c  �\   �M�f��U���U�E�E��}� t@�M����t6�E����E��M�;Mr�#  �U�E�f�f�
�U���U�E����E����M�M��}� t�U����t5�M����.t*�E����E��M�;Mr��   �.   �E�f��M���M�U����t6�M����M��U�;Ur�   �E�M�f�f��E���E�M����M����U����U��E�;Ev�e3ɋU�f�
�}�tP�}���tG�E�;Es?�M+M�9��s����U��	�E+E��E�M���Qh�   �U��E�PQ�S�����3���   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R�����������t3�t	�E�   ��E�    �U܉U�}� uh��j jlh�xj�&�������u̃}� u-����� "   j jlh�xh`xh���������"   ��   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�E�    �E�    �E�    �} u�e  �} u�} u�} t�} u�H  �} u�} u�} t�} u�+  �} u�}  u�} t�}  u�  �}$ u�}( u�}$ t�}( u��  �}� ��   �E�   �E�E�}� v�M����t�E���E�M���M��܋U����:u2�} t!�}s�  j�MQ�UR�EP��������M���M�_�} tY3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E؋M���Qh�   �U��R�������E�    �E�    �E�E��	�M���M�U����t4�M����/t�E����\u�U���U���E����.u�U�U�빃}� t>�} t0�E�+E���E��M;M�w�  �U�R�EP�MQ�UR��������E��E�_�} tY3ɋUf�
�}�tK�}���tB�}v<�E��9��s����M��	�U���UԋE���Ph�   �M��Q�������}� ty�U�;Urq�} t0�E�+E���E��M ;M�w��   �U�R�EP�M Q�UR�F������}$ t0�E�+E����E��M(;M�w�   �U�R�E�P�M(Q�U$R�������   �} t0�E�+E���E��M ;M�w�   �U�R�EP�M Q�UR��������}$ tX3��M$f��}(�tJ�}(���tA�}(v;�U(��9��s
����E��	�M(���MЋU���Rh�   �E$��P�������3��  �E�   �} t_�} vY3ɋUf�
�}�tK�}���tB�}v<�E��9��s����M��	�U���ŰE���Ph�   �M��Q臽�����} t_�} vY3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���EȋM���Qh�   �U��R�"������} t^�}  vX3��Mf��} �tJ�} ���tA�} v;�U ��9��s
����E��	�M ���MċU���Rh�   �E��P込�����}$ t_�}( vY3ɋU$f�
�}(�tK�}(���tB�}(v<�E(��9��s����M��	�U(���U��E���Ph�   �M$��Q�Y�����3҃} �U��}� u!h�yj h�   hhyj蠻������u̃}� u3�����    j h�   hhyhDyh�y�	������   �   �}� tw3�t	�E�   ��E�    �U��U܃}� u!hyj h�   hhyj� �������u̃}� u0�����    j h�   hhyhDyhy�������   ��Q���� "   �"   ��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�} t��}��E�P�V  ���M��} t
��  �U���]��������������������������̋�U�����}��E�P�
  ���E��=<� t�]�M�Q��  ��E���E���]�������������������������������̋�U��QV�}���=<� t�E�P�  �����w  ����M�Q�  ��^��]�������������������������������̋�U����} t^��}��E�P��  ���E�M#M�U��#U�ʉM��E�;E�t'�M�Q�Z  ��f�E��m���}��U�R�  ���E��E�M���} t)�=<� t�UR�EP��  ���M��	�U�    �   ��]��������������������������������������������̋�U��E%����P�MQ������]��������������������̋�U�����}��E�P��  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�`  ��f�E��m���}��U�R�  ���E�=<� tB�EP�MQ��  ���E�U�# z�E�# z;�t�E�E�   ����E�E����E��]������������������������������������������������̋�U����} 	 u>�}�u8��}��E�%=  ==  u$�=<� t�]��M�����  ���  u�;��7j h[  h�zh�zh(z�U������R�EPj �&�����P��������]��������������������������������������̋�U���荷��� �E����I����R	  �}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]�������������������������̋�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]��������������������������������������������������������������������������������������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��������������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�������������������������������������̋�U��Q�����E��E�P�)  ����]������������������̋�U��Q�]��e���U��E�P��  ����]��������������̋�U����E%�E�]��M�Q�   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R��  ���E��E�P�K������]��M�Q�2   ����]�������������������������������������������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]��������������������������������������������������������������������������������������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]��������������������������������������������������������������������������������������������̋�U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]��������������������������������������������̋�U��Q�E��  �E�P��������]�������������������̋�U��h4��EP�MQ�E�����]��������������������̋�U���<���3ŉE�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U܋E�H�M��U����E�}����u8�E�    �M�Q�x�������t	�E�    ��U�R�Z������E�   �Z  �E�P�M�Q�ǣ�����U�U؋E�HQ�U�R�W�������t	�E���E�M�U�A+B9E�}�M�Q��������E�    �E�   ��   �U�E�;Bk�M�Q�U�R�V������E؉E�M�Q+U�UċE�P�M�Q苺�����U�BP�M�Q�ʸ�����U�B��P�M�Q�b������E�    �E�   �~�U�E�;|B�M�Q�\������U܁�   ��U܋E�HQ�U�R�������E��UJ�M��E�   �2�E�M�H�M��U܁�����U܋E�HQ�U�R�۹�����E�    �E�H���    +щU��E��M���E܋M���Ɂ�   ���EԋU�z@u�E�MԉH�U�E����M�y u�U�Eԉ�E��M�3��"�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ��������u�U�R�EP�������E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������������������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]��������������������������������������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P�:������E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R��������E��ȋE���]������������������������������������������������������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]����������������̋�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]����������������������������������̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�����������������������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]������������������������������������������������������������������̋�U��hL��EP�MQ�������]��������������������̋�U������3ŉE��E�    �E�H
���  f�M��U�B
% �  f�E�M�Q�U�E�H�M�U����E�j@�M�Q�`�������t�E�   �f�U�f��f�U��E�=�  u�E�   �M�U�Q�E�M��U��E�ЋMf�Q�E��M�3��n�����]��������������������������������������������������������������̋�U���   ���3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!h0|j h�   h�{j��������u̃}� u0�J����    j h�   h�{hh{h0|�R�����3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$��.
�U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p������.
�$��.
�E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h�����/
�$�/
�E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d�����d/
�$�X/
�E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q�f������}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�|�����f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3�莓����]Ë�J&
�&
�'
)(
)
*
?*
$+
�*
w+
�,
 ,
�'
|'
�'
�'
  ��(
�(
�(
  ��)
�)
�)
  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U������3ŉE�����`�E��} u�   �} }�M�ىM�h���`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP誨����눋M�3��������]�����������������������������������������������������������̋�U���L���3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�f������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q茘����f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R�`�����f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3��ʊ����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]������������������������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]���������������������������̋�U������3ŉE��EPj j j �MQ�UR�EP�M�Q������ �E�UR�E�P�[������E��}�u	�M���M�E�M�3��V�����]��������������������������������������̋�U���x���3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|h�}h�}h�}ht}j�U��R觤����P�������E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   h�}h�}h }h}j�U��R�H�����P艖�����E�@�E�    �   �}�   �uK�}� uEj h�   h�}h�}h�|h�|j�M��Q������P�2������U�B�E�    �Cj h�   h�}h�}h`|hX|j�E��P謣����P�������M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q�'������U����?  |f�E�f��f�E��M�Q�U�R襞�����Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R�ː������}� },�E���%�   �E��	�M����M��}� ~�U�R赈������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P�V������M�Q�J������U�R�E�P�Q������M�Q�.������U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3�苂����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����EP�M�R�E�Q�׏�����E��}� t0�U��Rj�E�HQ趏�����E��}� t�U�B���M�A�U��R�E�HQ�U�BP聏�����E�}� t�M�Q���E�P�M��Q�U�BP�M�QR�L�������]�������������������������������������������������̋�U����֍����   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR�؇�����   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�i   �� �   ��]���������������������������������������������������������������������������������������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}��3����E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  膋�����    u��  �s������   �E�e������   �M�E�j�UR�׃������t�����E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u�P���������    ty�������   �E��؊��ǀ�       �M�Q�UR��  ������t�C�M�Q�  ���Ѕ�t+j�EP�^�����h�~�M��>���h���M�Q������x����U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP胑�����E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q蹐������u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�  ��,�	���D���������M��tj�UR誔�����E�����   �M��������!���   �E�x ��   �M�QR�EP��  ���ȅ���   荈�����   �U��������   �E��q����M���   �c����U���   �}$ u�EP�MQ荒����UR�E$P�~���j��MQ�UR�EP虂�����M�QR�C  �������M���   � ����U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP�  �� �軁��谇�����    u���{����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�M��EP�M��,����M���~�E���]� ��������̋�U��Q�M��E�� �~�M��
�����]������������������̋�U��Q�M��M��(����E��t�M�Q�*�����E���]� �����������������̋�U��Q�M��EP�M��p����M���~�E���]� ��������̋�U���V�E�8  �u�c  腅�����    tW�w������҂��9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP�U������t��   �M�y t��ly���U�R�E�P�MQ�U R�EP�w������E���M����M��U����U��E�;E���   �M��U;|\�E��M;HQ�U��B�����M��Q�| t�E��H�����U��B�L�Q��u�E��H�����U��B���@t�w���j�U$R�E P�M�Qj �U��B�����M�AP�UR�EP�MQ�UR�EP��  ��,�3���^��]���������������������������������������������������������������������������������������������������������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�[~������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����������������������������������������������������̋�U����E��M��U���E��}�RCC�t(�}�MOC�t�}�csm�t�@虂��ǀ�       �|��腂�����    ~�w����   �E�M����E�3��3���]�������������������������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E��ʁ���   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}���u���M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R��{���E�    ��E�P藊����Ëe��E�    �M��M��f����E������   �)�������    ~�����   �EԋUԋ���MԉËU�;Uu��%u���E�M�H�M�d�    Y_^[��]������������������������������������������������������������������������������������������������̋�U����E�E��}  t�M Q�UR�E�P�MQ袏�����}, u�UR�EP�Z�����MQ�U,R�K����E$�Q�UR�EP�M�Q�bz�����U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�T   ���E��}� t�EP�M�Q�s����]�������������������������������������������������������̋�U��j�h@�h9�d�    P���SVW���1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R�A}�����E���~�����   �E���~�����   �M���~���U���   ��~���M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP誉�����E��E�    ��   �M�Q�N  ��Ëe��u~��ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP�(x�����E�    �E�    �E������E�    �   �   �M�U��Q��E�P�\������q}���Mȉ��   �c}���Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP�b������t�M�Q�UR轈����ËEЋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u��{��ǀ     �   ��3���]�����������������������������������̋�U��j�hp�h9�d�    P���SVW���1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR�zs������t9j�E�P�Vv������t'�M��U�B��M��Q�U��P�o�����M����o���@  �U���txj�M�QR�s������tYj�E�P��u������tG�M�QR�E�HQ�U�R��z�����E�xu"�M��9 t�U��R�E��Q� o�����U����n���   �E�x uZj�M�QR�r������t>j�E�P�su������t,�M�QR�E��P�M�QR��n����P�E�P�Oz������n���[j�M�QR�=r������tAj�E�P�u������t/�M�QR�˂������t�E���t	�E�   ��E�   ��m���E�������   Ëe��Us���E������E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j�h��h9�d�    P���SVW���1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�������E��}�t�}�t+�R�U��R�E�HQ��l����P�U�BP�M�Q�|���)j�U��R�E�HQ�l����P�U�BP�M�Q�m���E�������   Ëe��q���E������M�d�    Y_^[��]��������������������������������������������������������������������̋�U��j�h��h9�d�    P��SVW���1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR�Jn���E�������E�����Ëe��p���E������M�d�    Y_^[��]�������������������������������������������������̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]������������������������̋�U����u��3Ƀ��    ����]������̋�U���(�} u3���  �E��M��} t�U�B����   �M��9MOC�t�U��:RCC�t�E��@uz�M��9csm�uK�U��zuB�E��x �t�M��y!�t�U��z"�u�E��x u�Mu�����    u3��I  �8u���   �E܋M܋���E܉�   �%  �M��9csm��  �U��z�  �E��x �t�M��y!�t�U��z"���   �E��x u#��t�����    u3���   �t�����   �M��U�U�E�E��M���   ��M��U��B�H���M�U��B�H��U���E����E��M���M�}� ~d�U��E��M��QR�E�P�M�Q�{������t?�2t���   �E؋U؋���M؉�} t�U�R�E�P�MQ�U�R�z������   ��3���]�����������������������������������������������������������������������������������������������������������������������������̋�U����E�    �E�E��M����M�U���U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u��r�����   �E��M��QR�E�P�q�����E���r���M􋐈   ��r���M����   ��r���M����   ��U�������E�� �����r���   �E�M����E��hr�����    }�Zr��ǀ�       �   ��]������������������������������������������������������������������������������������̋�U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!�q���   �E��U�����M���   �3���]����������������������������������������������̋�U����E�E��M����M�U���U��E�8��G  �M�Q��t�����} ��   ��p�����   �:csm�u~��p�����   �xum��p�����   �y �t(��p�����   �z!�t�p�����   �x"�u1�p�����   �QR��r������tj�p�����   P�:|�����kp�����   �9csm�um�Xp�����   �zu\�Gp�����   �x �t(�3p�����   �y!�t�p�����   �z"�u �} t�p���   �E��E�����U��
��o���M����   ��o���M�����   ��]���������������������������������������������������������������������������������������������������������̋�U��   ]����̋�U��j�hЬh9�d�    P��SVW���1E�3�P�E�d�    �e��E�    �M�U�E�������E�P�ix����Ëe��E������M�d�    Y_^[��]��������������������������������������������̋�U��j�h�h9�d�    P��SVW���1E�3�P�E�d�    �e��E�    �EP�U���E�������M�Q��w����Ëe��E������M�d�    Y_^[��]����������������������������������������̋�U��j�h�h9�d�    P��SVW���1E�3�P�E�d�    �e��E�    �EP�U�E�������M�Q�(w����Ëe��E������M�d�    Y_^[��]�������������������������������������������̋�U��j�h0�h9�d�    P��SVW���1E�3�P�E�d�    �e��E�    �EP�MQ�UR�EP�U�E�������M�Q�|v����Ëe��E������M�d�    Y_^[��]�����������������������������������������������̋�U����} t��a���} u�f���E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR�s������t�E���뀊E��]������������������������������������������������������������̋�U��j�h /d�    PQSVW���3�P�E�d�    �e��k�����    u���_���E�    ��g���$�k���M���   j j ��k���E������id
��E������[e���M�d�    Y_^[��]������������������������������������������������̋�U��Q�E�    �	�E����E��M�U�;}'hp��E����M�Q�L��w������t����2���]���������������������������������̋�U����} t���^���E��M�}� t���^���U�:csm�u/�E�xu&�M�y �t�U�z!�t�E�x"�u��^���M�Q�B���E��M�Q�B��M���U����U��E����E��}� ~0�M���U��E��H��Q�M��r��P��d������u�   ��3���]�����������������������������������������������������������U���SQ�E���E��EU�u�M�m���l��VW��_^��]�MU���   u�   Q�l��]Y[�� �������������������̋�U��=�� uj �EP�MQ�URhH��:   ����j �EP�MQ�URj �   ��]�������������������������̋�U��j�hX/d�    P��lVW���3�P�E�d�    �EP�M��.j���E�    �} t�M�U�3��} ���E��}� uhDwj j^h�~j�`������u̃}� uN�qw���    j j^h�~h�~hDw�|q�����E�    �E�    �E������M��w���E��U��<  �} t�}|�}$~	�E�    ��E�   �U��U��}� uhXvj j_h�~j�p_������u̃}� uN��v���    j j_h�~h�~hXv��p�����E�    �E�    �E������M��w���E��U��  �M�M��E�    �E�    �U���E�M����M��M��Z^����t0�M��N^������   ~�M��;^��Pj�E�P��q�����E��j�M�Q�M��^��P�qX�����E��}� t�U���E�M����M���U��-u�E���E�M���U�E����E���M��+u�U���E�M����M��} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E����E��M���U�E����E��E�RPj�j���s���E�U�j�M�Q�M��]��P�lW������t�U��0�U��Th  �E�P�M���\��P�AW������t0�M��a|�U��z�E�� �E���M�M��U���7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u^�U�;U�uV�u�3��E�RPj�j��}t���u��}��E��U��E�;E�w.r�M�;M�w$�E�RP�U�R�E�P�\���M�3��։EĉU���U���U�} u��E���M�U����U�������E����E��M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�zs��� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M���U��t�E��؋Mȃ� �ىEĉMȋUĉU��EȉE��E������M��~s���E��U��M�d�    Y_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�EP�t�����]���������������̋�U��=�� uj�EP�MQ�URhH��:�������j�EP�MQ�URj ������]�������������������������̋�U��j�EP�MQ�UR�EP�������]���������������̋�U��Q�E�    ��E����E��M���M�U�;Us�E���t�ڋE���]��������������������̋�U���<�EP�M���b���} u�E�    �M���p���E��  3Ƀ} ���M�}� uh�j j=hpj�X������u̃}� u=�
p���    j j=hphLh��j�����E�����M��fp���E��  3��} ���E�}� uh j j>hpj�6X������u̃}� u=�o���    j j>hphLh �i�����E�����M���o���E��!  ����;U����E�uh,j j?hpj��W������u̃}� u=�$o���    j j?hphLh,�/i�����E�����M��o���E��   �M���V���P�z u(�EP�MQ�UR�EP�T�����E̍M��Do���E��u�M��V���H�QR�EP�MQ�UR�EPh  �M��V���H�QR�M��wV��P�yX���� �E��}� u�E�����M���n���E���E����EčM���n���Eċ�]����������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�h����]�������������������̋�U����E�    � ��E��M��9 ��   j j j j j��U��Pj j ���E�}� u����   j=h�jj�M�Q�Gl�����E��}� u����rj j �U�R�E�Pj��M��Rj j ����uj�E�P�c��������=j �M�Q�Em������}�}� tj�U�R�nc�����E�    �E����E��4���3���]�����������������������������������������������������������������������̋�U��3�]��������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^����������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�����������������̋�U���(�E�E��M�M��U�U��}��g  �E��$�u
�M�Q�U�R��  ���E�}� t�E�E��s�M���Q�U���R��  ���E�}� t�E�E��F�M���Q�U���R�  ���E�}� t�E�E���M���Q�U���R�  ���E�E�E�M�M�E���   �U�R�E�P�Y  ���E�}� t�M�M��F�U���R�E���P�2  ���E�}� t�M�M���U���R�E���P�  ���E܋M܉M��E��i�U�R�E�P��   ���E�}� t�M�M���U���R�E���P��   ���E؋E��*�M�Q�U�R�   ���3���EP�M�Q�U�R�  ����]Ð�t
�t
�t
*t
�s
�����������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��+�P�   ����]�����������������̋�U��} t3��} ���D ��E�E]����������������̋�U����} �R  �EP�MQ�Q	  ���E��}� t�E��O  �U��R�E��P�*	  ���E��}� t�E��(  �M��Q�U��R�	  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�g  ���E��}� t�E��e  �U��R�E��P�@  ���E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$��|
�U��R�E��P��  ���E��}� t�E���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��}  �U��R�E��P�X  ���E��}� t�E��V  �M��Q�U��R�1  ���E��}� t�E��/  �E��P�M��Q�
  ���E��}� t�E��  �U��R�E��P��  ���E��}� t�E���  3���  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q�  ���E��}� t�E��  �U��R�E��P�g  ���E��}� t�E��e  �M��Q�U��R�@  ���E��}� t�E��>  �E��P�M��Q�  ���E��}� t�E��  �U��	R�E��	P��  ���E��}� t�E���  �M��Q�U��R��  ���E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R�b  ���E��}� t�E��`  �E��P�M��Q�;  ���E��}� t�E��9  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���E��}� t�E���  �E��
P�M��
Q��  ���E��}� t�E���  �U��R�E��P�  ���E��}� t�E��  �M��Q�U��R��  ���  �E��P�M��Q�]  ���E��}� t�E��[  �U��R�E��P�6  ���E��}� t�E��4  �M��Q�U��R�  ���E��}� t�E��  �E��P�M��Q��  ���E��}� t�E���   �U��R�E��P��  ���E��}� t�E��   �M��Q�U��R�  ���E��}� t�E��   �E��P�M��Q�s  ���E��}� t�E��t�U��R�E��P�o������E��}� t�M��M��F�U��R�E��P�H������E��}� t�M��M���U��R�E��P�!������E��M��M�E��3���]Ë��x
�y
�z
|
zx
�y
�z
�{
Sx
ky
�z
�{
,x
Dy
pz
�{
x
y
Iz
u{
�w
�x
"z
N{
�w
�x
�y
'{
�w
�x
�y
 {
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U���M��;�tK�E�E��M�M�U�R�E�P�������E�}� t�M�M���U���R�E��P�\������E�E��3���]�������������������������������������������̋�U��� �E�E��M�M��U��E��
;��   �U�U��E�E�M�Q�U�R��������E�}� t�E�E��s�M���Q�U��R�������E�}� t�E�E��F�M���Q�U��R�������E�}� t�E�E���M���Q�U��R�n������E��E��E�M�M�E��3���]�����������������������������������������������������������������̋�U����6O���   �E��} u�E�P�\  ���  �M��U��E��@�M��A�U��z t#�E��H���t�E���Pjhh���  ���M��A    �U��: ��   �E�������   �E��x t�M��Q���t�M�Q�O  ����U�R�	  ���E��x uG�M�Qj@h���u  ����t0�U��z t�E��H���t�E�P��  ����M�Q�1	  ���0�U��z t�E��H���t�E�P�  ����M�Q�?  ���U��z u3��N  �} t�E�   �E���E�    �M�Q�U�R�U  ���E��}� t!�}���  t�}���  t�E�P�4��u3���   j�M��QR����u3���   �} t&�E�M�f�Qf��E�M�f�Qf�P�Ef�M�f�H�} ��   �U�=  u4j h1  hЊh��hx�h\�j@�MQ�G]����P�O����� j@�URh  �E��HQ����u3��Bj@�U��@Rh  �E��HQ����u3��j
j�U�   R�E�P�:W�����   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�   �E�    �E�;Eb�}� t\�E�E�+����E��M��U��P�M�R�Z�����E�}� u�E��M�T��E���}� }�M����M�	�U����U��3��}� ����]�����������������������������������̋�U��Q�E�Q��E����3҃��E�P�M�QR��E����3Ƀ����U�J�E�@    �M�y t	�E�   ��U�P��  ���E��M�U��Qjhp�
���E�H��   t�U�B%   t�M�Q��u
�E�@    ��]����������������������������������������������������������̋�U���   ���3ŉE��9J���   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q����u��|����B    �   �  �E�P��|����QR�X�������r  jx�E�P��|����Q��ҁ������  R��x���P����u��|����A    �   �G  �U�R��|����Q�;X������u:��|����B  ��|����A��|�����x����B��|�����x����Q��   ��|����H����   ��|����z tt��|����HQ�U�R��|����Q�7O������uQ��|����B����|����A��|�����x����B��|����R�iC������|���;Au��|�����x����B�E��|����Q��u7��x���P��  ����t$��|����Q����|����P��|�����x����Q��|����H��   ��   ��  jx�U�R��|����H��Ɂ������  Q��x���R����u��|����@    �   �  �M�Q��|����P�V�������
  ��|����Q��   ��|����P��|����y t7��|����B   ��|����A��|����z u��|�����x����H�   ��|����z tl��|����Q�B������|���;BuP��|���Pj��x���Q��  ����t2��|����B   ��|����A��|����z u��|�����x����H�2��|����B   ��|����A��|����z u��|�����x����H�   ��|����z ut��|����x th�M�Q��|����P�oU������uO��|���Qj ��x���R�C  ����t3��|����H��   ��|����J��|����x u��|�����x����Q��|����@��������M�3��x8����]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�E�Q�?����3҃��E�P�M�y t	�E�   ��U�P��  ���E��M�U��Qjh`�
���E�H��u
�U�B    ��]��������������������������������������������̋�U���   ���3ŉE��ID���   ��|����EP�  ����x���jx�M�Q��|����B���%���  P��x���Q����u��|����B    �   �  �E�P��|����R�R������u`��|����x u��|���Qj��x���R�y  ����t3��|�����x����H��|�����x����B��|����Q����|����P�   ��|����y ut��|����z th�E�P��|����R� R������uO��|���Pj ��x���Q��  ����t3��|�����x����B��|�����x����Q��|����H����|����J��|����@��������M�3��)5����]� ������������������������������������������������������������������������������������������������������̋�U��E�HQ�=����3҃��E�Pjh��
���M�Q��u
�E�@    ]��������������������������̋�U���   ���3ŉE���A���   ��|����EP�B  ����x���jx�M�Q��|����B���%���  P��x���Q����u��|����B    �   �s�E�P��|����QR�SP������uF��x���P��  ����t3��|�����x����Q��|�����x����H��|����B����|����A��|����B��������M�3��e3����]� ������������������������������������������������������������������̋�U��Q�E�H��  �U�J�d�E��E�M��H�U�E��B��]�������������������������̋�U��Q�} t�E���thL��UR�E;������u0j�E�Ph  �M�QR����u3��Y�}� u�(�K�FhH��EP� ;������u"j�M�Qh   �U�BP����u3����MQ�oN�����E��E���]��������������������������������������������������������̋�U���f�Ef�E��E�    �	�M����M��}�
s�U��E��ED�;�u3���ظ   ��]����������������������̋�U���V�E%�  �ȁ�   �щU�j�E�Ph   �M�Q����u3��9�U;U�t,�} t&�E�Q��   �����U�P�9����;�u3���   ^��]������������������������������������̋�U����E�    �E��M��U��E���E��tM�M���a|�U���f�E���'�E���M���A|�U���F
�E����E��M����U��DЉE�뚋E���]������������������������������������̋�U����E�    �E��M��U���U�E���A|	�M���Z~�U���a|%�E���z�M����M��U��E��M���M���E���]�������������������������̋�U��Q���P�l�E��}� t�U�j��7����jj �>2�����4/����]�������������������̋�U��Q�E�    ���P�l�E��MQ������E���]��������������̋�U����P�l]�������������̋�U���   ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M���=���E�    �K���E�3Ƀ} �������������� u!h�j h  h��j��3������u̃����� uF�;K���    j h  h��hP�h��CE����ǅ8��������M��K����8����  3��} �������������� u!ht�j h  h��j�U3������u̃����� uF�J���    j h  h��hP�ht��D����ǅ4��������M��	K����4����z  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���h  ������ �[  �������� |%��������x�������� ���� ����
ǅ ���    �� ���������������k�	�������� ����������������   3�tǅ���   �
ǅ���    ����������������� u!h j ha  h��j��1������u̃����� uF�EI���    j ha  h��hP�h �MC����ǅ0��������M��I����0����  �����������������*  ������$���
�E�   ������Q�UR������P�Y  ����  �E�    �MЉMԋUԉU�E�E��E�    �E������E�    ��  ������������������ ����������wL�������4�
�$��
�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��M  ��������*u(�UR�E�����E�}� }�E����E��M��ىM���U�k�
�������LЉM��   �E�    ��  ��������*u�EP�fE�����Ẽ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  �������\�
�$�H�
�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��v
  ������������������A����������7�J  �������Ȥ
�$���
�M���0  u	�U��� �U��E�   �EP�C����f�������M��� tW���������   ������ƅ���� �M��-��P�M��-��� ���   Q������R������P��C������}�E�   �f������f�������������U��E�   �  �EP�C���������������� t�������y u� ��U��E�P�0�����E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�Ủ�����������|����MQ�7B�����E��U��� ��   �}� u� ��E��M��������E�    �	�U܃��U܋E�;�|���}L���������t?�M��,��P�������Q��-������t������������������������������d�}� u	���M��E�   �U���x�����|�����|�������|�����t��x������t��x�������x����ɋ�x���+U����U��  �EP�1A������t����O8������   3�tǅ���   �
ǅ���    �������p�����p��� u!h�j h�  h��j�+������u̃�p��� uF��B���    j h�  h��hP�h���<����ǅ,��������M��MC����,����  ��  �M��� t��t���f������f����t�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}̣   ~Ah�  h��j�Ḿ�]  Q�f$�����E��}� t�U��U��E�]  �E���Ẹ   �M���M�U�B��J���h�����l����M��)��P�U�R�E�P������Q�U�R�E�P��h���Q�H�R�l�Ѓ��E�%�   t%�}� u�M��W)��P�M�Q�T�R�l�Ѓ���������gu)�M���   u�M��!)��P�U�R�P�P�l�Ѓ��M����-u�E�   �E��M����M��U�R�,�����E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�/������X�����\����   �U���   t�EP��.������X�����\����   �M��� tB�U���@t�EP�=��������X�����\�����MQ�=���������X�����\����=�U���@t�EP�n=�������X�����\�����MQ�S=����3҉�X�����\����E���@t@��\��� 7|	��X��� s,��X����ً�\����� �ډ�P�����T����E�   �E����X�����P�����\�����T����E�% �  u&�M���   u��P�����T����� ��P�����T����}� }	�E�   ��M�����M��}�   ~�E�   ��P����T���u�E�    �������E��M̋Ũ��U̅���P����T���t{�E��RP��T���Q��P���R�>����0��d����E��RP��T���P��P���Q�=����P�����T�����d���9~��d����������d����E���d�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅L����M���u������R�EP��L���Qj �N  ���U�R������P�MQ�U�R�E�P�  ���M���t$�U���u������P�MQ��L���Rj0�  ���}� ��   �}� ��   �E���H����M܉�D�����D�����D�������D�����~}�M��$��P�M��$������   R��H���P������Q��:������@�����@��� ǅ���������2������R�EP������Q��  ����H����@�����H����j�����E�P������Q�UR�E�P�M�Q�v  �������� |$�U���t������P�MQ��L���Rj ��  ���}� tj�E�P�2�����E�    �s��������� t������tǅ ���    �
ǅ ���   �� �����<�����<��� u!h�j h�  h��j��#������u̃�<��� uC�P;���    j h�  h��hP�h��X5����ǅ(��������M��;����(������������$����M��;����$����M�3��$����]��
/�
b�
ؖ
%�
1�
t�
��
��
��
��
��
ʖ
Ӗ
 �I �
��
��
��
��
 �i�
�
2�
/�
��
��
 �
�
r�
v�
(�
E�
�
;�
"�
   	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ��/�����Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U����E�    �E�    �E�H��pt	�U��pu�E�H�U3�;����#  �E�H��st�U�B��St	�E�    ��E�   �M�M��U��st�E��St	�E�    ��E�   �M��M��}� u�}� tA�U�;U�u*�E�H�� ��Ƀ��U�� ��҃�;�u	�E�   ��E�    �E��  �E�H��dtv�U�B��itj�M�Q��ot^�E�H��utR�U�B��xtF�M�Q��Xt:�E��dt1�M��it(�U��ot�E��ut�M��xt�U��X��   �E�H��dtE�U�B��it9�M�Q��ot-�E�H��ut!�U�B��xt�M�Q��Xt	�E�    ��E�   �E��dt6�M��it-�U��ot$�E��ut�M��xt�U��Xt	�E�    ��E�   �E�;E�t3��T�M�Q��   ����ڋE%   �����;�u�M�Q�� ����ڋE�� �����;�t3���M�3�;U����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����  ���3ŉE�ǅ4���    ǅ����    ǅ����    ǅd���    ǅ����    ǅl���    ǅ����    �EP��T����"��ǅ����    ǅt���    ǅ@���    ǅ����    ǅx�������ǅ��������ǅ��������ǅp�������ǅ��������ǅ����    ��/����|���3Ƀ} ����0�����0��� u!h�j h  h��j�(������u̃�0��� uI�/���    j h  h��hp�h��)����ǅ,���������T�����/����,����3  3��} ����,�����,��� u!ht�j h  h��j�������u̃�,��� uI��.���    j h  h��hp�ht��)����ǅ(���������T����N/����(����3  ǅL���    �U������ǅ@���    ���@�������@�����@�����2  ��@���u������ u�2  ǅ����    ǅ8���    ǅ����    ǅP���    ǅx�������ǅ����    ǅd���    �������Mǅ��������ǅ��������ǅp�������ǅ���������Uf�f��D�����D����U���U���K/  ��L��� �>/  ��D����� |%��D�����x��D����� ���������
ǅ����    ��������H�����H���k�	��8����� ����8�����8�����  �U���%��  �������u\j
��t���Q�UR�������~9��t������$u+��@��� uh@  j ������R�����ǅ����   �
ǅ����    �������)  j
��t���P�MQ�F��������������t������U��@��� ��   ������ |#��t������$u������d}ǅ����   �
ǅ����    ��������(�����(��� u!h(!j hQ  h��j�������u̃�(��� uI�,���    j hQ  h��hp�h(!�&����ǅ$���������T����i,����$����40  ������;�x���~���������������x�����������������x����   ��8�����   3�tǅ����   �
ǅ����    ��������$�����$��� u!h j h]  h��j��������u̃�$��� uI�.+���    j h]  h��hp�h �6%����ǅ ���������T����+���� ����L/  ��8����������������N,  �������$�X�
��@��� u	������t��@���u�������u�,  ǅ����   ��L���Q�UR��D���P�=  ����+  ǅh���    ��h�����l�����l���������������������ǅ����    ǅd�������ǅ����    �+  ��D����������������� ������������wj����������
�$�x�
���������������E���������������4���������������#�������ʀ   ����������������������	+  ��D�����*��  ������ u�UR�0'�����������`  j
��t���P�MQ����������������t������U��@��� ��  ������ |#��t������$u������d}ǅ|���   �
ǅ|���    ��|����� ����� ��� u!hp j h�  h��j�M������u̃� ��� uI�(���    j h�  h��hp�hp �"����ǅ���������T�����(���������,  ������;�x���~��������x������x�����x�����x�����x����������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R���������؉����u!h�j h�  h��j�������u̃���� uI�r'���    j h�  h��hp�h��z!����ǅ���������T�����'��������+  �(  �+������������������������P��$���������������� }���������������������ډ������������k�
��D����TЉ������2(  ǅd���    �#(  ��D�����*��  ������ u�MQ�J$������d����`  j
��t���R�EP����������p�����t������M��@��� ��  ��p��� |#��t������$u������d}ǅt���   �
ǅt���    ��t������������� u!hj h�  h��j�g������u̃���� uI��%���    j h�  h��hp�h������ǅ���������T����&���������)  ��p���;�x���~��p�����p������x�����p�����p�����x�����p����������� uG��p�����Ǆ����   ��p�����f��D���f��������p������������������   ������Q��D���Rj��p�����������Q�0��������؉����u!hhj h�  h��j�.������u̃���� uI�$���    j h�  h��hp�hh�����ǅ���������T�����$��������(  ��%  �+��p���������������������R��!������d�����d��� }
ǅd����������d���k�
��D����TЉ�d����_%  ��D�����l�����l�����I��l�����l���.�D  ��l�������
�$���
�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������d�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu������   �������ǅ8���    ������#�������� ���������������   ��������#  ��D�����h�����h�����A��h�����h���7�B!  ��h�����$�
�$���
��������0  u�������� ������ǅ����   ������ u�EP������f��<�����  ������ |������d}ǅd���   �
ǅd���    ��d������������� u!hj hv  h��j�!
������u̃���� uI�!���    j hv  h��hp�h�����ǅ���������T�����!��������%  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P���������؉����u!h�j hz  h��j�	������u̃���� uI�m ���    j hz  h��hp�h��u����ǅ���������T����� ��������$  �  �,���������������� ����� ���Q������f��<����������� t_��<���%�   ������ƅ���� ��T�������P��T����������   R������P��P���Q�������}
ǅl���   �f��<���f��P�����P���������ǅ����   �^  ������ u�MQ�������������  ������ |������d}ǅ`���   �
ǅ`���    ��`��������������� u!hj h�  h��j�y������u̃����� uI�����    j h�  h��hp�h������ǅ���������T����*���������"  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�i��������؉�����u!h j h�  h��j�g������u̃����� uI�����    j h�  h��hp�h ������ǅ ���������T�������� �����!  �w  �+��������������������������R����������������� t�������x u#� �������������R������������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q��������������������  ��������0  u�������� ��������d����uǅ\���������d�����\�����\��������������� u�EP�������������  ������ |������d}ǅX���   �
ǅX���    ��X��������������� u!hj h6  h��j�z������u̃����� uI�����    j h6  h��hp�h������ǅ����������T����+����������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�j��������؉�����u!h j h:  h��j�h������u̃����� uI�����    j h:  h��hp�h ������ǅ����������T��������������  �x  �+��������������������������Q������������������� ��   ������ u� �������������������ǅ����    ���������������������;�����}O���������tB��T�������P�������Q�������t������������������������������v������ u��������ǅ����   ����������������������������������t���������t���������������ɋ�����+��������������'  ������ u�EP��������������  ������ |������d}ǅT���   �
ǅT���    ��T��������������� u!hj h�  h��j�B������u̃����� uI����    j h�  h��hp�h�����ǅ����������T��������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�2	��������؉�����u!h j h�  h��j�0 ������u̃����� uI����    j h�  h��hp�h �����ǅ����������T��������������  �@  �+��������������������������Q�������������������   3�tǅP���   �
ǅP���    ��P��������������� u!h�j h�  h��j�O�������u̃����� uI����    j h�  h��hp�h������ǅ����������T���� ����������  �_  �������� t������f��L���f����������L����ǅl���   �%  ǅh���   ��D����� f��D�����������@��������������  ��@��� ��  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u!hj h�  h��j��������u̃����� uI�z���    j h�  h��hp�h�����ǅ����������T��������������  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������R��D���Pj��������������R���������؉�����u!hxj h�  h��j��������u̃����� uI�u���    j h�  h��hp�hx�}����ǅ����������T��������������  �'  ��P���������ǅP���   ��d��� }ǅd���   �7��d��� u��D�����guǅd���   ���d���   ~
ǅd���   ��d����   ~Yh�  h��j��d���]  P������������������ t ��������������d�����]  ��P����
ǅd����   ������ u#�E���E�M�Q��A��������������  ������ |������d}ǅH���   �
ǅH���    ��H��������������� u!hj h  h��j�o�������u̃����� uI�����    j h  h��hp�h������ǅ����������T���� ����������  ��@���t!h8j h  h��j���������u̋����������������������������������������Q��A���������������T�������P��h���Q��d���R��D���P��P���Q������R������P�H�Q�l�Ѓ���������   t.��d��� u%��T�������P������P�T�Q�l�Ѓ���D�����gu2������%�   u%��T����x���P������Q�P�R�l�Ѓ����������-u!��������   ��������������������������Q��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅd���   ǅ4���   �
ǅ4���'   ǅ����   ������%�   t&�0   f��������4�����Qf������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  �%  ������ u�EP��������������������  ������ |������d}ǅD���   �
ǅD���    ��D��������������� u!hj h�  h��j�_�������u̃����� uI����    j h�  h��hp�h��	����ǅ����������T��������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�O ��������؉�����u!h�j h�  h��j�M�������u̃����� uI����    j h�  h��hp�h������ǅ����������T���������������  �]  �1��������������������������Q�������������������  ��������   �%  ������ u�EP���������������������  ������ |������d}ǅ@���   �
ǅ@���    ��@��������������� u!hj h�  h��j�(�������u̃����� uI����    j h�  h��hp�h�����ǅ����������T��������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P����������؉�|���u!h�j h�  h��j��������u̃�|��� uI�t���    j h�  h��hp�h��|����ǅ����������T��������������  �&  �1����������������x�����x���Q���������������������  �������� �e  ��������@�)  ������ u�MQ�	��������������������  ������ |������d}ǅ<���   �
ǅ<���    ��<�����t�����t��� u!hj h�  h��j���������u̃�t��� uI�A���    j h�  h��hp�h�I����ǅ����������T�������������_  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�����������؉�p���u!h�j h�  h��j���������u̃�p��� uI�/
���    j h�  h��hp�h��7����ǅ����������T����
���������M  ��  �3����������������l�����l���R��������������������(  ������ u!�EP�`���������������������  ������ |������d}ǅ8���   �
ǅ8���    ��8�����h�����h��� u!hj h�  h��j��������u̃�h��� uI�	���    j h�  h��hp�h�����ǅ����������T����i	���������4  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P����������؉�d���u!h�j h�  h��j��������u̃�d��� uI����    j h�  h��hp�h������ǅ����������T����W���������"  �  �5����������������`�����`���Q�]��������������������Z  ��������@�'  ������ u�EP�$�������������������  ������ |������d}ǅ4���   �
ǅ4���    ��4�����\�����\��� u!hj h  h��j��������u̃�\��� uI�����    j h  h��hp�h�� ����ǅ����������T����0����������
  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������P��D���Qj��������������P�o���������؉�X���u!h�j h  h��j�m�������u̃�X��� uI�����    j h  h��hp�h��������ǅ����������T��������������	  �}  �2����������������T�����T���Q�$������������������$  ������ u�UR������3ɉ�������������  ������ |������d}ǅ0���   �
ǅ0���    ��0�����P�����P��� u!hj h0  h��j�W�������u̃�P��� uI����    j h0  h��hp�h������ǅ����������T��������������  ��@��� �  �������������� uG��������Ǆ����   ��������f��D���f���������������������������   ������Q��D���Rj��������������Q�G���������؉�L���u!h�j h4  h��j�E�������u̃�L��� uI����    j h4  h��hp�h�������ǅ����������T���������������  �U  �3����������������H�����H���R�� ����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ��������������d��� }ǅd���   �%�����������������d���   ~
ǅd���   �����������u
ǅ����    ��O�����������d�����d�������d������������������   �������RP������P������Q�����0�������������RP������R������P�v ��������������������9~�������4�������������������������������������K�����O���+���������������������������������   t>������ t���������0t'���������������������0��������������������u��@��� u�k  ��l��� �:  ��������@tj��������   t�-   f������ǅ����   �D��������t�+   f������ǅ����   �!��������t�    f������ǅ����   ������+�����+�������D�����������u��L���Q�UR��D���Pj ��  ����|���Q��L���R�EP������Q������R�  ����������t'��������u��L���R�EP��D���Qj0�  �������� ��   ������ ��   ��������@�����������<�����<�����<�������<�������   ��T����x���P��T����l���� ���   Q��@���R��<���P���������8�����8��� ǅL��������2��L���Q�UR��<���P�E  ����@����8�����@����`����(��|���R��L���P�MQ������R������P��  ����L��� |'��������t��L���R�EP��D���Qj �T  �������� tj������R�S�����ǅ����    ������8��� t��8���tǅ,���    �
ǅ,���   ��,�����4�����4��� u!h�j h�  h��j��������u̃�4��� uI�����    j h�  h��hp�h�������ǅ����������T����e����������0  �������  ��@��� ��  ǅ����    ���������������������;�x�����  ����������������(�����(�������(�����(�����   ��(����$�\�
���������E�������MQ��������_  ���������E�������MQ��������;  ���������E�������MQ�������  ���������E�������MQ��������   ���������E�������MQ�b�������   ���������E�������MQ��������������������   3�tǅ$���   �
ǅ$���    ��$�����0�����0��� u!hpj h.	  h��j��������u̃�0��� uF�����    j h.	  h��hp�hp������ǅ����������T����Y����������'�����#�����L�����������T����0����������M�3��������]Ë�"�
u�
ƴ
Z�
1�
@�
�
v�
!�
2�
�
��
F�
U�
 �I }�
N�
A�
_�
q�
 ���
��
8�
�
��
��
м
��
��
\�
��
U�
��
�
��
   	
��
��
��

�
.�
��
R�
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�H��@t�U�z u�E����U�
�4�EP�MQ�7������Ё���  u�E� ������M����E�]����������������������������������̋�U��E�M���M��~!�UR�EP�MQ�Y������U�:�u���]������������������������̋�U����E��M��U�B��@t�M�y u�U�E�M��y�U�    �E�M���M��~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������렋E�8 u�M�U����]������������������������������������������������̋�U��j�h�h9�d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� uh8�j j3h��j�X�������u̃}� u-�����    j j3h��h��h8�����������  �M�U�U�E�P�\������E�    �M�Q�UR������f�E��E������   ��E�P�I������f�E��M�d�    Y_^[��]����������������������������������������������������������������������������̋�U���8���3ŉE�V�E�H��@�d  �UR�`��������t@�EP�O��������t/�MQ�>����������UR�-�������������E���E���E�H$�����у�tj�EP����������t@�MQ����������t/�UR������������EP���������������E���E���M�Q$������uh�M�Q���U��E�M��H�}� |2�U�f�Mf��U����  f�UދE����U�
f�E��  ��EP�MQ��������  �(  �UR�$��������t@�EP���������t/�MQ�����������UR���������������E���Eب��E��H��   ��   �URj�E�P�M�Q��������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���UԋE�MԉH�}� |.�U��M��T��E�����   �UЋE����U�
��EP�M��T�R�������EЃ}��u���  �k�|����E%��  �[�E�H���M̋U�ẺB�}� |/�M�f�Ef��M����  f�MʋU����M�f�E����UR�EP�:�����^�M�3��0�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EP�MQ�c�����]��������̋�U��j j jj jh   @h��`���]����������̋�U��=���t�=���t���P��]������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��������������������������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]������������������̋�U����E��t
�-���]���M��t����-���]������U��t
�-���]���E��t	�������؛�M�� t���]����]�������������������������̋�U��Q�=<� t�]���E�    �E���]�������������̋�U��j�h �h9�d�    P���SVW���1E�3�P�E�d�    �e�=<� ��   �E��@tp�=�� tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe����    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]�������������������������������������������������������̋�U��Q�=<� t�]��e���U���]�����������������̋�U��Q�=<� t�����E��E���?�E���E�    �E���]����������������̋�U��Q�=<� t������E��E���?�E�������E�    �E���]���������������������������̋�U����=<� t8�����E��E#E�M��#M���E��U������U��U��E�P�e�������E�    �E���]�������������������������̋�U��Q�����E��E��?E��E��M�Q��������]����������������������̋�U������3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ�������UR�������E�P�MQ�������UR�������E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR� �����f�E�f��f�E��؋Mf�U�f�Q
�M�3��n�����]����������������������������������������������������������������������������������������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��� VW�   �(��}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q�_^��]� ���������������������̋�U��Q�M��E�� T��M��A    �U��B �E���]����������������������̋�U��Q�M��M��C����E��t�M�Q�������E���]� �����������������̋�U��Q�M��E�� T��M��A    �U��B �E�Q�M�������E���]� ���������������������̋�U��Q�M��E�� T��M��U��A�M��A �E���]� ������������������̋�U��Q�M��E�� T��M��A    �U��B �EP�M��M����E���]� �����������������������̋�U��Q�M��E�;Et0�M������M�Q��t�E�HQ�M��������U��E�H�J�E���]� ���������������������̋�U��Q�M��E�� T��M��3�����]������������������̋�U����M��E��x t�M��Q�U���E�`��E���]�������������������̋�U����M��} tK�EP�(��������E��M�Q�������U��B�E��x t�MQ�U�R�E��HQ�g������U��B��]� �����������������������������̋�U��Q�M��E��H��t�U��BP�4������M��A    �U��B ��]������������������������̋�U��Q�M��EP�M��l����M��|��E���]� ��������̋�U��Q�M��M������E��t�M�Q�������E���]� �����������������̋�U��Q�M��EP�M�������M��|��E���]� ��������̋�U��Q�M��E�� |��M��������]������������������̋�U��Q�M��EP�M������M�����E���]� ��������̋�U��Q�M��M��g����E��t�M�Q��������E���]� �����������������̋�U��Q�M��EP�M������M�����E���]� ��������̋�U��Q�M��E�� ���M��
�����]������������������̋�U��Q�M��EP�M��<����M�����E���]� ��������̋�U��Q�M��M��?����E��t�M�Q��������E���]� �����������������̋�U��Q�M��EP�M�������M�����E���]� ��������̋�U��Q�M��E�� ���M�������]������������������̋�U����EP�M������M$Q�U R�EP�MQ�UR�EP�MQ�M��-���P�2   �� �E�M������E��]�����������������������������̋�U���8���3ŉE�} ~�EP�MQ�K  ���E��}�}3��<  �}  ~�U R�EP�#  ���E ��} �}3��  �E�    �}$ u�M��B�E$�} t
�}  �j  �M;M u
�   ��  �} ~
�   ��  �}~
�   �  �U�R�E$P�0��u3��  �} u�} t-�}u�}  t!h�j h�   h��j�|�������u̃} ~m�}�s
�   �R  �U։U��	�E���E�M����t8�E��H��t-�U��M��;�|�E��U��B;�
�   �  뵸   ��  �}  ~m�}�s
�   ��  �M։M��	�U���U�E����t8�U��B��t-�M��E��;�|�U��M��Q;�
�   �  뵸   �  j j �EP�MQj	�U$R��E��}� u3��Z  �}� ~63�u2�����3��u���r#h��  �M��T	R�P�����P�w������E���E�    �ẺE��}� u3��  �M�Q�U�R�EP�MQj�U$R���u
��   ��   j j �E P�MQj	�U$R��E�}� u
�   �   �}� ~63�u2�����3��u��r#h��  �M�T	R������P��������E���E�    �EȉE��}� u�O�M�M�Q�U�R�E P�MQj�U$R���t!�E�P�M�Q�U�R�E�P�MQ�UR�\�E�E�P�*������M�Q�������E�M�3�謸����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]��������������������������̋�U���<�EP�M������} u�E�    �M������E��  3Ƀ} ���M�}� uhp�j j?h��j�Y�������u̃}� u=�����    j j?h��hԍhp���������E�����M������E��  3��} ���E�}� uh��j j@h��j��������u̃}� u=�G����    j j@h��hԍh���R������E�����M������E��.  ����;U����E�uh�uj jAh��j�s�������u̃}� u=������    j jAh��hԍh�u��������E�����M��0����E��   �M�蓺����z u-�M�胺��P�EP�MQ�UR�ܳ�����E̍M�������E��~�M��V���� �HQ�UR�EP�MQ�URh  �M��3���� �HQ�M��%���P�'����� �E��}� u�����    �E�����M������E���U����UčM��p����Eċ�]�������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��=�� u�EP�MQ�UR�X�������j �EP�MQ�UR������]������������������̋�U���$V�E�    �E�    3��} ���E܃}� uh̐j jThX�j�C�������u̃}� u.�����    j jThX�h<�h̐����������T  �U��E�}� tj=�M�Q�ÿ�����E��}� t�U�;U�u�I����    ����  �E�+E�=�  |h��j jfhX�j褸������u�h�  �U���R������=�  rh��j jghX�j�k�������u̋M��Q��҃��U���;��u���Q�g  ������=�� ��   �} t*�= � t!�f�����t�{����    ����F  �   �}� t3��4  �   �=�� u8h�   hX�jj貱��������=�� u�����  ����    �= � u7h�   hX�jj�q������ ��= � u����  � ��     ����M��}� u-3�u!h �j h�   hX�j�5�������u̃���r  �M�+M�Q�U�R�  ���E�}� ��   �E��8 ��   j�M�U���P�������}� ti�	�M���M�U�E��<� t�M�U��E�u��D����ց}����?s2h�   hX�jj�M�Q���R�������E��}� t�E������M�U��E���M�    �   �}� ��   �}� }�U��ډU�E��;E�|:�M�������?s,h�   hX�j�U��Rj���P螮�����E��}� u����D  �M�U��E���M�U��D�    �E�     �M�����j�U�R��������E�     3���   �} ��   h  hX�jj�M�Q蚸������P�%������E�}� ��   j h  hX�h<�h���U�R�E�P�[�������P�M�Q�������P�������U�+U�U�U��E��  �M����M��U������#U�R�E�P����u�E������}��u�[���� *   j�M�Q�������}� tj�U�R��������E�     �E�^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q����E��	�M����M��U��: tK�EP�M��R�EP�3�������u/�M���E���=t�U���M���u�E�+�����뤋E�+�����؋�]����������������������������������̋�U����E�    �E�E�} u3���   �M��E���E��t�M����M���h�  hX�jj�U���R� ������E��E��E��}� u
j	��������M�M�U�: ��   �E�Q�P��������E�h�  hX�jj�U�R��������M���U��: t7j h�  hX�hd�h���E�Q�U�R�E��Q�l�����P譼�����U���U�E����E��k����M��    �E���]��������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�   ��]�������������������̋�U���$�} t�E�M�3҃} �U�}� uhDwj j^h��j���������u̃}� u-�U����    j j^h��h��hDw�`�����3��'  �} t�}|�}$~	�E�    ��E�   �M��M�}� uhXvj j_h��j�u�������u̃}� u-������    j j_h��h��hXv�������3��  �E�E��E�    �M�f�f�U��E����E�j�M�Q螺������t�U�f�f�E��M����M����U���-u�E���E�M�f�f�U��E����E���M���+u�U�f�f�E��M����M��} u@�U�R�"�������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q�ܭ������u2�U����xt�M����Xu�E����E��M�f�f�U��E����E����3��u�E��M�Q莭�����E��}��t�V�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��E܋M܃�7�M���h�U�;Ur�^�E���E�M�;M�r�U�;U�u���3��u9U�w�E��EE��E���M���M�} u��U�f�f�E��M����M��*����U����U��E��u�} t�M�M��E�    �f�U��u*�E��uV�M��t	�}�   �w�U��u=�}����v4�V���� "   �E��t	�E�������M��t	�E�   ���E�����} t�U�E���M��t�U��ډU�E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�UR�X�����]�������������������̋�U��j�EP�MQ�UR�(�����]�������������������̋�U��j�EP�MQ�UR�������]�������������������̋�U��� �} uh`�j jdhX�j��������u̋M�M��U�R�������E��E��H��   u&�2���� 	   �U��B�� �M��A���  �c  �/�U��B��@t$����� "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�`����� 9E�t�S�����@9E�u�M�Q��������u�U�R詸�����E��H��  �  �U��E��
+Hy!h��j h�   hX�j�i�������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P輩�����E��s�}��t!�}��t�M����U���������U���E���E��H�� t9jj j �U�R�������E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q�������E�U�;U�t�E��H�� �U��J���  ��E%��  ��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���0�EP�M��O���3Ƀ} ���M�}� uh��j j:h(�j�F�������u̃}� u=觿���    j j:h(�h�h��貹�����E�    �M������E���   �M��f����@�x u#�MQ�UR�8������E��M��Ͽ���E���   �	�E���E�Mf�f�U��E���t|�M������H�U��D��tS�M���M�U���u�E�    �M��n����E��j�M����U��9Mu�M���M؍M��D����E��@��U�9Uu��h����E�9Eu�M�MԍM������E���E�    �M������EЋ�]���������������������������������������������������������������������������������������������������������̋�U��j �EP�MQ�i�����]�������̋�U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[������������������������������������������������������%h�%l�%p�%t�%x�%|�%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��% �%�%�%�%�%�%�%�% �%$�%(�%,�%0�%4�%8�%<�%@�%D�%H�%L�%P�%T�%X�%\�%`�%d�%h�%l�%p�%t�%x�%|�%��%��%��%��%��%��%��%��%��%��%��%��%d�%`�%\�%������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍M������T$�B�J�3�賓��� ��J���������������̍M������T$�B�J�3�胓��� �����������������̡��������ËT$�B�J�3��M����Ъ��������������������������̍M��z����T$�B�J�3��������骫��������������̋T$�B�J�3��������邫����������������������̍M������T$�B�J�3�賒������J������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������p��H�_^[��]����������������U����   SVW��@����0   �������x��0�_^[��]����������������U����   SVW��@����0   ����������@�_^[��]����������������U����   SVW��@����0   ����������8�_^[��]����������������U����   SVW��@����0   ����������X�_^[��]����������������U����   SVW��@����0   ����������P�_^[��]����������������U����   SVW��@����0   ����������(�_^[��]����������������U����   SVW��@����0   ��������� �_^[��]����������������U����   SVW��@����0   ������� ����_^[��]����������������U����   SVW��@����0   �������(����_^[��]����������������U����   SVW��@����0   �������H����_^[��]����������������U����   SVW��@����0   �������P����_^[��]����������������U����   SVW��@����0   �������h����_^[��]����������������U����   SVW��@����0   �������p����_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ����������x�_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   �����������_^[��]����������������U����   SVW��@����0   ������� ����_^[��]����������������U����   SVW��@����0   �������8�� �_^[��]����������������U����   SVW��@����0   �������@����_^[��]����������������U����   SVW��@����0   �������`����_^[��]����������������U����   SVW��@����0   �������h����_^[��]����������������U����   SVW��@����0   �������P��@�_^[��]����������������U����   SVW��@����0   �������X��(�_^[��]����������������U����   SVW��@����0   �������x��8�_^[��]����������������U����   SVW��@����0   ����������0�_^[��]����������������U����   SVW��@����0   ����������P�_^[��]����������������U����   SVW��@����0   ����������H�_^[��]����������������U����   SVW��@����0   ���������� �_^[��]����������������U����   SVW��@����0   �������ȅ��_^[��]����������������U����   SVW��@����0   ������� ����_^[��]����������������U����   SVW��@����0   ���������x�_^[��]����������������U����   SVW��@����0   �������(����_^[��]����������������U����   SVW��@����0   �������0����_^[��]����������������U����   SVW��@����0   �������H����_^[��]����������������U����   SVW��@����0   �������P����_^[��]����������������U����   SVW��@����0   �������p��p�_^[��]����������������U����   SVW��@����0   �������x��h�_^[��]����������������U����   SVW��@����0   �������h����_^[��]����������������U����   SVW��@����0   �������p����_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   �������؇���_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   �������`��@�_^[��]����������������U����   SVW��@����0   �������h���_^[��]����������������U����   SVW��@����0   ����������0�_^[��]����������������U����   SVW��@����0   ���������� �_^[��]����������������U����   SVW��@����0   ����������P�_^[��]����������������U����   SVW��@����0   ����������H�_^[��]����������������U����   SVW��@����0   �������Ј��_^[��]����������������U����   SVW��@����0   �������؈��_^[��]����������������U����   SVW��@����0   ������h    jjj��v����P��v����P��v�����8�_^[���   ;��9�����]�������������������������������������U����   SVW��@����0   �������~���(�_^[���   ;��ه����]���������������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ����������x�_^[��]����������������U����   SVW��@����0   �������ȉ���_^[��]����������������U����   SVW��@����0   �������Љ���_^[��]����������������U����   SVW��@����0   �����������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ���������p�_^[��]����������������U����   SVW��@����0   ���������h�_^[��]����������������U����   SVW��@����0   �������X����_^[��]����������������U����   SVW��@����0   �������`����_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   �������Ȋ���_^[��]����������������U����   SVW��@����0   �������Њ���_^[��]����������������U����   SVW��@����0   ���������8�_^[��]����������������U����   SVW��@����0   ��������� �_^[��]����������������U����   SVW��@����0   �������0��0�_^[��]����������������U����   SVW��@����0   �������8��(�_^[��]����������������U����   SVW��@����0   �������P��H�_^[��]����������������U����   SVW��@����0   �������X��@�_^[��]����������������U����   SVW��@����0   �������x���_^[��]����������������U����   SVW��@����0   �����������_^[��]����������������U����   SVW��@����0   ����������p�_^[��]����������������U����   SVW��@����0   ����������X�_^[��]����������������U����   SVW��@����0   ����������h�_^[��]����������������U����   SVW��@����0   ���������`�_^[��]����������������U����   SVW��@����0   ������� ����_^[��]����������������U����   SVW��@����0   ���������x�_^[��]����������������U����   SVW��@����0   �������(��P�_^[��]����������������U����   SVW��@����0   �������0��H�_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ����������p�_^[��]����������������U����   SVW��@����0   ������������_^[��]����������������U����   SVW��@����0   ���������x�_^[��]����������������U����   SVW��@����0   ������� ����_^[��]����������������U����   SVW��@����0   �����������_^[��]����������������U����   SVW��@����0   �������(��h�_^[��]����������������U����   SVW��@����0   �������0��`�_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �?�?@P@�@�@APA        �A�ABPB�B�BCPC        �C�CDPD�D�DEPE        �E�EFPF�F�FGPG        �G�GHPH�H�HIPI        �I�IJPJ�J�JKPK        �K�KLPL�L�LMPM�MN        `N�N�N O`O�O�O P        `P�P�P Q`Q�Q�Q R        `R�R�R S`S�S�S T        `T�T�T U`U�U�U V        `V�V�V W`W�W�W X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��'�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ����                                                                                                                                                                                                                                                                    Z�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ���R       X   ܗ ��                                                                                                                                                                              	              	            	              	         ?             @                  �   &   ��������5            4  �������5            4  �������                                                 	       ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                       �        �������                        ��������       ����    ���� �  �      ��� �         �        �������                        ��������       ����    ���� �  �      ��� �  Can't load anima dlls       .cdl    Anima.C4D15     \   found programPath %s
       PATH    Anima.xml File not found!
      Anima.xml File not found!       an(i)ma StartupError        r   Anima.xml   c4d_main        ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                      �?                        ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                c:\lavoro\anima\sdk\src\resource\_api\c4d_basebitmap.cpp            Stop    Stop:   res c:\lavoro\anima\sdk\src\resource\_api\c4d_misc\datastructures\basearray.h               ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                            c:\lavoro\anima\sdk\src\resource\_api\c4d_file.cpp              Debug Stop      Debug Stop:         c:\lavoro\anima\sdk\src\resource\_api\c4d_misc\memory\defaultallocator.h                ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                               %s  c:\lavoro\anima\sdk\src\resource\_api\c4d_general.h                 ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                            
   CRITICAL:       WARNING:     [%s %s L%d]    %H:%M:%S    c:\lavoro\anima\sdk\src\resource\_api\c4d_misc\memory\debugglobals.cpp                  ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                            H��    ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                                ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                            c:\lavoro\anima\sdk\src\resource\_api\c4d_string.cpp            no baselist         ����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?                            f c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c                       ( s t r e a m   ! =   N U L L )         _ f c l o s e _ n o l o c k         ( s t r   ! =   N U L L )               (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       (   s t r   ! =   N U L L   )           (   c o u n t   > =   0   )         f g e t s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f g e t s . c                     (   s t r i n g   ! =   N U L L   )   | |   (   c o u n t   = =   0   )                 ( * m o d e   ! =   _ T ( ' \ 0 ' ) )           ( m o d e   ! =   N U L L )         _ f s o p e n       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f o p e n . c                     ( f i l e   ! =   N U L L )         f o p e n _ s       ( p f i l e   ! =   N U L L )           p r i n t f     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ p r i n t f . c                       ( f o r m a t   ! =   N U L L )             f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c                            �    s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y [ n ] )                       s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y _ a b b r [ n ] )                         _ G e t d a y s _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r f t i m e . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\strftime.c               s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h [ n ] )                     s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h _ a b b r [ n ] )                       _ G e t m o n t h s _ l             s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w w _ t i m e f m t )                     s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w w _ l d a t e f m t )                           s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w w _ s d a t e f m t )                           s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > a m p m [ 1 ] )                   s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > a m p m [ 0 ] )                   s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > m o n t h [ n ] )                         s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > m o n t h _ a b b r [ n ] )                       s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w d a y [ n ] )                   s t r c p y _ s ( s ,   l e n   -   ( s   -   p ) ,   p t - > w d a y _ a b b r [ n ] )                     _ G e t t n a m e s _ l         F A L S E           ( " I n v a l i d   M B C S   c h a r a c t e r   s e q u e n c e   p a s s e d   t o   s t r f t i m e " , 0 )                         t i m e p t r   ! =   N U L L           (   f o r m a t   ! =   N U L L   )             (   m a x s i z e   ! =   0   )         _ S t r f t i m e _ l       (   s t r i n g   ! =   N U L L   )                 (   " I n v a l i d   f o r m a t   d i r e c t i v e "   ,   0   )                     (   t i m e p t r - > t m _ y e a r   > =   - 1 9 0 0   )   & &   (   t i m e p t r - > t m _ y e a r   < =   8 0 9 9   )                           (   t i m e p t r - > t m _ y e a r   > = 0   )             (   (   t i m e p t r - > t m _ s e c   > = 0   )   & &   (   t i m e p t r - > t m _ s e c   < =   5 9   )   )                         (   (   t i m e p t r - > t m _ m i n   > = 0   )   & &   (   t i m e p t r - > t m _ m i n   < =   5 9   )   )                         (   (   t i m e p t r - > t m _ y d a y   > = 0   )   & &   (   t i m e p t r - > t m _ y d a y   < =   3 6 5   )   )                           (   (   t i m e p t r - > t m _ h o u r   > = 0   )   & &   (   t i m e p t r - > t m _ h o u r   < =   2 3   )   )                             (   (   t i m e p t r - > t m _ m d a y   > = 1   )   & &   (   t i m e p t r - > t m _ m d a y   < =   3 1   )   )                             (   (   t i m e p t r - > t m _ m o n   > = 0   )   & &   (   t i m e p t r - > t m _ m o n   < =   1 1   )   )                         _ e x p a n d t i m e           (   (   t i m e p t r - > t m _ w d a y   > = 0   )   & &   (   t i m e p t r - > t m _ w d a y   < =   6   )   )                               ( " I n v a l i d   M B C S   c h a r a c t e r   s e q u e n c e   p a s s e d   i n t o   s t r f t i m e " , 0 )                             ( " I n v a l i d   M B C S   c h a r a c t e r   s e q u e n c e   f o u n d   i n   l o c a l e   A M P M   s t r i n g " , 0 )                               a/p am/pm       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h                           ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                   _ g e t _ t i m e z o n e ( & t i m e z o n e )             _ g e t _ d s t b i a s ( & d s t b i a s )             _ g e t _ d a y l i g h t ( & d a y l i g h t )             (   p t i m e   ! =   N U L L   )           _ l o c a l t i m e 6 4 _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c t i m 6 4 . c                       (   p t m   ! =   N U L L   )           ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                 _ v s n p r i n t f _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c                       ����    f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c          _ g e t _ e r r n o         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d o s m a p . c                       p V a l u e   ! =   N U L L         _ g e t _ d o s e r r n o           . . .       A s s e r t i o n   F a i l e d         E r r o r       W a r n i n g       (���    f:\dd\vctools\crt_bld\self_x86\crt\src\dbgrpt.c             ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       p f n N e w H o o k   ! =   N U L L             _ C r t S e t R e p o r t H o o k W 2               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c                           m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y                     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   ( * _ e r r n o ( ) )           D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )                                     
 M o d u l e :         
 F i l e :         
 L i n e :         
 
     E x p r e s s i o n :               
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                     m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                 < p r o g r a m   n a m e   u n k n o w n >                 w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       _ _ c r t M e s s a g e W i n d o w W           Client  Ignore  CRT Normal  Free    X�P�L�D�<�    Error: memory allocation: bad memory block type.
           Invalid allocation size: %Iu bytes.
        Client hook allocation failure.
        Client hook allocation failure at file %hs line %d.
            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c                         _ C r t C h e c k M e m o r y ( )           _ p F i r s t B l o c k   = =   p O l d B l o c k               _ p L a s t B l o c k   = =   p O l d B l o c k             f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       Error: possible heap corruption at or near 0x%p                 p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Client hook re-allocation failure.
         Client hook re-allocation failure at file %hs line %d.
             _ e x p a n d _ d b g       p U s e r D a t a   ! =   N U L L           _ p F i r s t B l o c k   = =   p H e a d           _ p L a s t B l o c k   = =   p H e a d             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                                 HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()                _ m s i z e _ d b g         %hs located at 0x%p is %Iu bytes long.
             %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
                   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 DAMAGED     _heapchk fails with unknown return value!
          _heapchk fails with _HEAPBADPTR.
       _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADBEGIN.
         _ C r t S e t D b g F l a g             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t D o F o r A l l C l i e n t O b j e c t s               p f n   ! =   N U L L       Bad memory block found at 0x%p.
        Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              _ C r t M e m C h e c k p o i n t           s t a t e   ! =   N U L L           n e w S t a t e   ! =   N U L L         o l d S t a t e   ! =   N U L L         _ C r t M e m D i f f e r e n c e           Object dump complete.
      crt block at 0x%p, subtype %x, %Iu bytes long.
             normal block at 0x%p, %Iu bytes long.
          client block at 0x%p, subtype %x, %Iu bytes long.
              {%ld}   %hs(%d) :       #File Error#(%d) :      Dumping objects ->
      Data: <%s> %s
     _ p r i n t M e m B l o c k D a t a             %.2X    Detected memory leaks!
     Total allocations: %Id bytes.
          Largest number used: %Id bytes.
        %Id bytes in %Id %hs Blocks.
       _ C r t M e m D u m p S t a t i s t i c s           o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g               Damage before 0x%p which was allocated by aligned routine
              The block at 0x%p was not allocated by _aligned routines, use realloc()                 The block at 0x%p was not allocated by _aligned routines, use free()                _ a l i g n e d _ m s i z e _ d b g             m e m b l o c k   ! =   N U L L             ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   ( _ o s f i l e ( f h )   &   F O P E N )           _ c l o s e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c                     ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     _ f i l e n o           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c                           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c                       s t r e a m   ! =   N U L L         _ f i l b u f       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f i l b u f . c                         s t r   ! =   N U L L       f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c             ccs UTF-8   UTF-16LE    UNICODE         ( * m o d e   = =   _ T ( ' \ 0 ' ) )           _ o p e n f i l e       ( " I n v a l i d   f i l e   o p e n   m o d e " , 0 )                 m o d e   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ o p e n . c                     f i l e n a m e   ! =   N U L L         f:\dd\vctools\crt_bld\self_x86\crt\src\stream.c             f:\dd\vctools\crt_bld\self_x86\crt\src\_sftbuf.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ s f t b u f . c                         f l a g   = =   0   | |   f l a g   = =   1             ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx                          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c             ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 ( c h   ! =   _ T ( ' \ 0 ' ) )         _ o u t p u t _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c                       v p r i n t f _ h e l p e r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v p r i n t f . c                         �h�    f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c           FlsFree     FlsSetValue     FlsGetValue     FlsAlloc    K E R N E L 3 2 . D L L         CorExitProcess      m s c o r e e . d l l       _ w p g m p t r   ! =   N U L L         _ g e t _ w p g m p t r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 d a t . c                         _ p g m p t r   ! =   N U L L           _ g e t _ p g m p t r       s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               _ s e t e n v p             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c                         f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c            f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c            f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c          f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h e a p i n i t . c                       _ c r t h e a p           �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �                                      Unknown Runtime Check Error
       Stack memory around _alloca was corrupted
         A local variable was used before it was initialized
           Stack memory was corrupted
            A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                x� �������`�                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                  Run-Time Check Failure #%d - %s         Unknown Module Name     Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s                   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                           Stack corrupted near unknown variable               Stack area around _alloca memory reserved by this function is corrupted
                %s%s%s%s    >   %s%s%p%s%ld%s%d%s       Stack area around _alloca memory reserved by this function is corrupted                 
Address: 0x    
Size:      
Allocation number within this function:            
Data: <    wsprintfA   u s e r 3 2 . d l l         A variable is being used without being initialized.             Stack around _alloca corrupted          Local variable used before initialization           Stack memory corruption     Cast to smaller type causing loss of data           Stack pointer corruption        ������d�<�    f:\dd\vctools\crt_bld\self_x86\crt\prebuild\misc\i386\chkesp.c                  The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                       _ s e t d e f a u l t p r e c i s i o n                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c                         s i z e I n B y t e s   >   0           _ c f t o e _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c                         b u f   ! =   N U L L       e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                           _ c f t o e 2 _ l           s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o a _ l         _ c f t o f _ l         _ c f t o f 2 _ l       _ c f t o g _ l         ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               B u f f e r   i s   t o o   s m a l l           ( ( ( _ S r c ) ) )   ! =   N U L L             s t r c p y _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l                           ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                     f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c            f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c a l r e f . c                       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )                                                                                         H H : m m : s s         d d d d ,   M M M M   d d ,   y y y y           M M / d d / y y         P M     A M     D e c e m b e r         N o v e m b e r         O c t o b e r       S e p t e m b e r       A u g u s t     J u l y     J u n e     A p r i l       M a r c h       F e b r u a r y         J a n u a r y       D e c       N o v       O c t       S e p       A u g       J u l       J u n       M a y       A p r       M a r       F e b       J a n       S a t u r d a y         F r i d a y     T h u r s d a y         W e d n e s d a y       T u e s d a y       M o n d a y     S u n d a y     S a t       F r i       T h u       W e d       T u e       M o n       S u n       HH:mm:ss    dddd, MMMM dd, yyyy     MM/dd/yy    PM  AM  December    November    October     September   August  July    June    April   March   February    January     Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday     Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec                _ g e t _ d a y l i g h t               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t i m e s e t . c                         ( _ D a y l i g h t   ! =   N U L L )           _ g e t _ d s t b i a s         ( _ D a y l i g h t _ s a v i n g s _ b i a s   ! =   N U L L )                 _ g e t _ t i m e z o n e           ( _ T i m e z o n e   ! =   N U L L )           _ I n d e x   = =   0   | |   _ I n d e x   = =   1             _ R e t u r n V a l u e   ! =   N U L L             _ g e t _ t z n a m e           ( _ B u f f e r   ! =   N U L L   & &   _ S i z e I n B y t e s   >   0 )   | |   ( _ B u f f e r   = =   N U L L   & &   _ S i z e I n B y t e s   = =   0 )                                   s t r n c p y _ s ( t z n a m e [ 1 ] ,   6 4 ,   T Z ,   3 )                   s t r n c p y _ s ( t z n a m e [ 0 ] ,   6 4 ,   T Z ,   3 )                   s t r c p y _ s ( l a s t T Z ,   s t r l e n ( T Z )   +   1 ,   T Z )                 f:\dd\vctools\crt_bld\self_x86\crt\src\tzset.c          TZ  _ t z s e t _ n o l o c k           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t z s e t . c                     _ i s i n d s t _ n o l o c k           c v t d a t e       s r c   ! =   N U L L       _ s t r i c m p _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r i c m p . c                         d s t   ! =   N U L L       _ s t r i c m p         (   t i m p   ! =   N U L L   )         _ g m t i m e 6 4 _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g m t i m e 6 4 . c                       _ g m t i m e 3 2 _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g m t i m e . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\gmtime.c             ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p                             p N o d e - > _ N e x t   ! =   N U L L                 s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ M _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                 f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c          f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t M o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c                         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   _ C r t S e t R e p o r t F i l e               _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                           s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 %s(%d) : %s         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed!       Assertion failed:       _CrtDbgReport: String too long or IO Error          s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   , Line      <file unknown>      Second Chance Assertion Failed: File            _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t A           w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               _CrtDbgReport: String too long or Invalid characters in String                  s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                       % s ( % d )   :   % s       w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                 w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d !           A s s e r t i o n   f a i l e d :                   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 
   ,   L i n e         < f i l e   u n k n o w n >             S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   _ V C r t D b g R e p o r t W           s i g n a l     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c                       ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f:\dd\vctools\crt_bld\self_x86\crt\src\winsig.c             r a i s e       GetProcessWindowStation     GetUserObjectInformationW       GetLastActivePopup      GetActiveWindow     MessageBoxW     U S E R 3 2 . D L L         ( s t r i n g   ! =   N U L L )         _ s w p r i n t f       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s w p r i n t f . c                       s i z e I n B y t e s   > =   c o u n t             m e m c p y _ s             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c                       w c s c p y _ s         ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ h a n d l e r . c p p                         p n h   = =   0         ... Assertion Failed    Error   Warning     ���    _ C r t S e t R e p o r t H o o k 2             Microsoft Visual C++ Debug Library              Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)                    
Module:    
File:      
Line:      

  Expression:     

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.                          <program name unknown>      s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         _ _ c r t M e s s a g e W i n d o w A           _ e x p a n d _ b a s e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c                       p B l o c k   ! =   N U L L         s p r i n t f           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s p r i n t f . c                         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c                         ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6             f:\dd\vctools\crt_bld\self_x86\crt\src\osfinfo.c            _ g e t _ o s f h a n d l e             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c                         ( _ o s f i l e ( f i l e d e s )   &   F O P E N )             _ c o m m i t           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c                           ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c                     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )               ( ( c n t   &   1 )   = =   0 )         _ w r i t e _ n o l o c k           ( b u f   ! =   N U L L )           ( c n t   < =   I N T _ M A X )         _ r e a d           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r e a d . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\read.c           ( i n p u t b u f   ! =   N U L L )             _ r e a d _ n o l o c k         f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c                         _ o p e n       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o p e n . c                       ( p a t h   ! =   N U L L )             ( ( p m o d e   &   ( ~ ( _ S _ I R E A D   |   _ S _ I W R I T E ) ) )   = =   0 )                     _ s o p e n _ h e l p e r           ( p f h   ! =   N U L L )           0   & &   " O n l y   U T F - 1 6   l i t t l e   e n d i a n   &   U T F - 8   i s   s u p p o r t e d   f o r   r e a d s "                               0   & &   " I n t e r n a l   E r r o r "           ( o f l a g   &   ( _ O _ T E X T   |   _ O _ W T E X T   |   _ O _ U 1 6 T E X T   |   _ O _ U 8 T E X T )   )   ! =   0                           (   " I n v a l i d   s h a r i n g   f l a g "   ,   0   )                 (   " I n v a l i d   o p e n   f l a g "   ,   0   )               _ g e t _ f m o d e ( & f m o d e )             _ t s o p e n _ n o l o c k         s 2   ! =   N U L L         _ m b s n b i c m p _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s n b i c m . c                       s 1   ! =   N U L L         _ m b s n b c m p _ l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s n b c m p . c                       _ i s a t t y           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c                       ( " B u f f e r   t o o   s m a l l " ,   0 )               _ w c t o m b _ s _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c                       s i z e I n B y t e s   < =   I N T _ M A X                 ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                           ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                   _ o u t p u t _ s _ l       ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 _ o u t p u t _ p _ l       f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c             r u n t i m e   e r r o r            
     T L O S S   e r r o r  
           S I N G   e r r o r  
         D O M A I N   e r r o r  
             R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                            �+   p+	    +
   �*   8*   �)   x)   )   �(   0(   �'   0'   �&   �&   �%    %!   �"x   �"y   �"z   \"�   T"�   0"                                        M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )                             w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )                                   w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )                           w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                             R u n t i m e   E r r o r ! 
 
 P r o g r a m :                     w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                     _ N M S G _ W R I T E           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c                         SystemFunction036       ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       A D V A P I 3 2 . D L L         r a n d _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ r a n d _ s . c                       _ R a n d o m V a l u e   ! =   N U L L             s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         _ _ g e t l o c a l e i n f o               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t h e l p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\inithelp.c           M S P D B 1 0 0 . D L L     M S V C R 1 0 0 D . d l l               PDBOpenValidate5    E n v i r o n m e n t D i r e c t o r y             S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 0 . 0 \ S e t u p \ V S                       RegCloseKey     RegQueryValueExW    RegOpenKeyExW   D L L       M S P D B 1 0 0         _ c o n t r o l f p _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c                           ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             p f l t   ! =   N U L L         s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           _ f p t o s t r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c                       s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                     _ f l t o u t 2             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c                         _ s e t _ o u t p u t _ f o r m a t             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t f o r m a t . c                               ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t t i m e . c                       p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                   f:\dd\vctools\crt_bld\self_x86\crt\src\inittime.c           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t n u m . c                         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initnum.c                f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t m o n . c                         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0               f:\dd\vctools\crt_bld\self_x86\crt\src\initmon.c                                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                            s t r n c p y _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l                         ( _ t c s n l e n ( o p t i o n ,   _ M A X _ E N V )   <   _ M A X _ E N V )                   g e t e n v     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t e n v . c                       ( o p t i o n   ! =   N U L L )             _ t c s n l e n ( * s e a r c h   +   l e n g t h   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                           s t r c p y _ s ( b u f f e r ,   s i z e I n T C h a r s ,   s t r )                   ( b u f f e r   ! =   N U L L   & &   s i z e I n T C h a r s   >   0 )   | |   ( b u f f e r   = =   N U L L   & &   s i z e I n T C h a r s   = =   0 )                                   _ g e t e n v _ s _ h e l p e r         p R e t u r n V a l u e   ! =   N U L L             s t r c p y _ s ( * p B u f f e r ,   s i z e ,   s t r )               v a r n a m e   ! =   N U L L           _ d u p e n v _ s _ h e l p e r         p B u f f e r   ! =   N U L L           p l o c i - > c t y p e 1 _ r e f c o u n t   >   0             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n i t c t y p . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\initctyp.c           LC_TIME     LC_NUMERIC      LC_MONETARY     LC_CTYPE    LC_COLLATE      LC_ALL      <L    �,L���� L����L��� L��Q��K����                	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         _ c o n f i g t h r e a d l o c a l e           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t l o c a l . c                       ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                       f:\dd\vctools\crt_bld\self_x86\crt\src\setlocal.c           s e t l o c a l e       L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     s t r n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ s e t l o c a l e _ n o l o c k           ;   =;  s t r c p y _ s ( p c h   +   s i z e o f ( i n t ) ,   c c h   -   s i z e o f ( i n t ) ,   l c t e m p )                         _ s e t l o c a l e _ s e t _ c a t             s t r c a t _ s ( p c h ,   c c h ,   " ; " )               _ s e t l o c a l e _ g e t _ a l l             =       s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   s t r n c p y _ s ( c a c h e i n ,   c a c h e i n S i z e ,   s o u r c e ,   c h a r a c t e r s I n S o u r c e   +   1 )                               C   s t r c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   " C " )                 _ e x p a n d l o c a l e           s t r c a t _ s ( o u t s t r ,   s i z e I n B y t e s ,   (   * ( c h a r   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( c h a r   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                           _ s t r c a t s             s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                               s t r n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   l o c a l e ,   l e n )                                             s t r n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   l o c a l e ,   l e n )                                           _., s t r n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & l o c a l e [ 1 ] ,   1 6 - 1 )                                             _ _ l c _ s t r t o l c         .   _   s t r c p y _ s ( l o c a l e ,   s i z e I n B y t e s ,   ( c h a r   * ) n a m e s - > s z L a n g u a g e )                         _ _ l c _ l c t o s t r         _ l s e e k i 6 4       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c                        Complete Object Locator'        Class Hierarchy Descriptor'         Base Class Array'       Base Class Descriptor at (          Type Descriptor'       `local static thread guard'         `managed vector copy constructor iterator'          `vector vbase copy constructor iterator'            `vector copy constructor iterator'          `dynamic atexit destructor for '        `dynamic initializer for '      `eh vector vbase copy constructor iterator'         `eh vector copy constructor iterator'           `managed vector destructor iterator'        `managed vector constructor iterator'           `placement delete[] closure'        `placement delete closure'      `omni callsig'       delete[]    new[]  `local vftable constructor closure'         `local vftable'     `RTTI   `EH `udt returning'     `copy constructor closure'      `eh vector vbase constructor iterator'          `eh vector destructor iterator'         `eh vector constructor iterator'        `virtual displacement map'      `vector vbase constructor iterator'         `vector destructor iterator'        `vector constructor iterator'       `scalar deleting destructor'        `default constructor closure'       `vector deleting destructor'        `vbase destructor'      `string'    `local static guard'        `typeof'    `vcall'     `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete      new    __unaligned     __restrict      __ptr64     __eabi  __clrcall   __fastcall      __thiscall      __stdcall   __pascal    __cdecl     __based(    �_�_�_�_�_�_�_�_�_�_x_k�p_d_ Q`_\_X_T_P_L_@_<_8_4_0_,_(_$_ ________ _�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^x^l^T^0^^�]�]�]t]T],]]�\�\�\�\�\�\T\L\@\,\\�[�[�[\[([[�Z�Z�ZLZ(Zk�Z�Y�Y�Y�Y                                                                                CV:     ::  '   `   generic-type-   template-parameter-     ''  `anonymous namespace'       `non-type-template-parameter        `template-parameter     void    NULL    extern "C"      [thunk]:    public:     protected:      private:    virtual     static      `template static data member destructor helper'             `template static data member constructor helper'            `local static destructor helper'        `adjustor{      `vtordisp{      `vtordispex{        }'  }'  )   void    std::nullptr_t      volatile    ,<ellipsis>     ,...    <ellipsis>       throw(      volatile   const   signed      unsigned    UNKNOWN     __w64   wchar_t     <unknown>   __int128    __int64     __int32     __int16     __int8  bool    double  long    float   long    int short   char    enum    cointerface     coclass     class   struct      union   `unknown ecsu'      int     short   char    const   volatile    cli::pin_ptr<   cli::array<     )[  {flat}  s   {for    ������    2�i�p�    ������    ���-�    H���*�     ??     ������    _ m b s t o w c s _ l _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c                       s   ! =   N U L L       r e t s i z e   < =   s i z e I n W o r d s             b u f f e r S i z e   < =   I N T _ M A X           _ m b s t o w c s _ s _ l           ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                                   ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               s t r c a t _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l                       _ v s n p r i n t f _ h e l p e r           s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   _ v s p r i n t f _ s _ l           f o r m a t   ! =   N U L L         _ v s n p r i n t f _ s _ l         l e n g t h   <   s i z e I n T C h a r s           2   < =   r a d i x   & &   r a d i x   < =   3 6                   s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   s i z e I n T C h a r s   >   0         x t o a _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c                       x 6 4 t o a _ s         _ w c s t o m b s _ l _ h e l p e r             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c                       p w c s   ! =   N U L L         s i z e I n B y t e s   >   r e t s i z e           _ w c s t o m b s _ s _ l           ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               w c s c a t _ s         _ v s w p r i n t f _ h e l p e r               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c                       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s w p r i n t f _ s _ l         _ v s n w p r i n t f _ s _ l           x t o w _ s     x 6 4 t o w _ s         _ w o u t p u t _ l         _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r             GetUserObjectInformationA       MessageBoxA     _ v s p r i n t f _ l       _ v s c p r i n t f _ h e l p e r               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c                           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                             ( s i z e   > =   0 )       _ c h s i z e _ s       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c h s i z e . c                       _ l s e e k         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k . c                     ( " I n v a l i d   f i l e   d e s c r i p t o r " , 0 )               _ s e t m o d e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t m o d e . c                         ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T )   | |   ( m o d e   = =   _ O _ U 8 T E X T )   | |   ( m o d e   = =   _ O _ U 1 6 T E X T ) )                                               _ s e t _ f m o d e         ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T ) )                             _ g e t _ f m o d e         ( p M o d e   ! =   N U L L )           c o u n t   < =   I N T _ M A X         _ s t r n i c m p _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c m p . c                       _ s t r n i c m p       i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                   s t r t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o l . c                       n p t r   ! =   N U L L         _ s e t _ e r r o r _ m o d e               f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c                         ( " I n v a l i d   e r r o r _ m o d e " ,   0 )               w c s n c p y _ s       _ w m a k e p a t h _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t m a k e p a t h _ s . i n l                         ( L " I n v a l i d   p a r a m e t e r " ,   0 )               _ w s p l i t p a t h _ s           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t s p l i t p a t h _ s . i n l                           ( ( ( _ P a t h ) ) )   ! =   N U L L                _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                         _ s e t _ c o n t r o l f p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                             _ _ s t r g t o l d 1 2 _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l                             _ L o c a l e   ! =   N U L L           1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 $ I 1 0 _ O U T P U T       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c                             ��bad exception   ������    s t r t o x q       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r t o q . c                       n   < =   I N T _ M A X         _ m b s n b i c o l l _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s n b i c o . c                       f:\dd\vctools\crt_bld\self_x86\crt\src\wtombenv.c           united-states   united-kingdom      trinidad & tobago       south-korea     south-africa    south korea     south africa    slovak  puerto-rico     pr-china    pr china    nz  new-zealand     hong-kong   holland     great britain   england     czech   china   britain     america     usa us  uk  swiss   swedish-finland     spanish-venezuela       spanish-uruguay     spanish-puerto rico     spanish-peru    spanish-paraguay    spanish-panama      spanish-nicaragua       spanish-modern      spanish-mexican     spanish-honduras    spanish-guatemala       spanish-el salvador     spanish-ecuador     spanish-dominican republic      spanish-costa rica      spanish-colombia    spanish-chile   spanish-bolivia     spanish-argentina       portuguese-brazilian        norwegian-nynorsk       norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg       german-lichtenstein     german-austrian     french-swiss    french-luxembourg       french-canadian     french-belgian      english-usa     english-us      english-uk      english-trinidad y tobago       english-south africa        english-nz      english-jamaica     english-ire     english-caribbean       english-can     english-belize      english-aus     english-american    dutch-belgian   chinese-traditional     chinese-singapore       chinese-simplified      chinese-hongkong    chinese     chi chh canadian    belgian     australian      american-english    american english    american    �ENU ؅ENU ąENU ��ENA ��NLB ��ENC ��ZHH ��ZHI ��CHS t�ZHH \�CHS D�ZHI ,�CHT �NLB �ENU ��ENA �ENL ԄENC ��ENB ��ENI ��ENJ ��ENZ l�ENS L�ENT <�ENG ,�ENU �ENU �FRB �FRC ܃FRL ̃FRS ��DEA ��DEC ��DEL x�DES h�ENI X�ITS L�NOR 8�NOR  �NON �PTB �ESS ؂ESB ȂESL ��ESO ��ESC |�ESD h�ESF P�ESE 8�ESG $�ESH �ESM ��ESN �ESI ЁESA ��ESZ ��ESR ��ESU ��ESY h�ESV T�SVF L�DES H�ENG D�ENU @�ENU                                                                                                         4�USA (�GBR  �CHN �CZE �GBR ��GBR ��NLD �HKG ԀNZL ЀNZL ĀCHN ��CHN ��PRI ��SVK ��ZAF ��KOR p�ZAF `�KOR H�TTO H�GBR 4�GBR $�USA D�USA                                     6-    Norwegian-Nynorsk           s t r c p y _ s ( l p O u t S t r - > s z L a n g u a g e ,   ( s i z e o f ( l p O u t S t r - > s z L a n g u a g e )   /   s i z e o f ( l p O u t S t r - > s z L a n g u a g e [ 0 ] ) ) ,   " N o r w e g i a n - N y n o r s k " )                                                   _ _ g e t _ q u a l i f i e d _ l o c a l e                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ g e t q l o c . c                         OCP ACP _ w o u t p u t _ s _ l         _ w o u t p u t _ p _ l         f p u t w c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f p u t w c . c                       C O N O U T $       csm�               �                ��0���    Unknown exception       ������    �o���    d�����    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ a _ c m p . c                     c c h C o u n t 1 = = 0   & &   c c h C o u n t 2 = = 1   | |   c c h C o u n t 1 = = 1   & &   c c h C o u n t 2 = = 0                             _ s t r i n g 2   ! =   N U L L         _ s t r n i c o l l _ l             f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t r n i c o l . c                       _ s t r i n g 1   ! =   N U L L         s t r c p y _ s ( n a m e ,   s t r l e n ( o p t i o n )   +   2 ,   o p t i o n )                     ( " C R T   L o g i c   e r r o r   d u r i n g   s e t e n v " , 0 )                   f:\dd\vctools\crt_bld\self_x86\crt\src\setenv.c                 _ t c s n l e n ( e q u a l   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                     e q u a l   -   o p t i o n   <   _ M A X _ E N V               _ _ c r t s e t e n v       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s e t e n v . c                       p o p t i o n   ! =   N U L L               s t r c p y _ s ( * n e w e n v p t r ,   e n v p t r S i z e ,   * o l d e n v p t r )                     c o p y _ e n v i r o n         w c s t o x l       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o l . c                       _ m b s c h r _ l           f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s c h r . c                       s t r i n g   ! =   N U L L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     RSDSe��,?�IJ�o˖�`O   C:\Lavoro\anima\sdk\src\Anima.Plugin\C4D\Debug\AnimaWrapper.pdb                                                                                                                                                                                                                                                                                                 p�`�               t�    |�    p�        ����    @   `�                    ����               ̙    ԙ    ��        ����    @   ��                    p��               $�    0�T�    p�       ����    @   �        ��        ����    @   x�                   ��    T�                ��x�                P�Ě               ؚ    �T�    P�       ����    @   Ě                    p� �               4�    @�T�    p�       ����    @    �                    ��|�               ��    ��@�T�    ��       ����    @   |�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ����    ����    ����    qK    ����    ����    ����    ZR    ����    ����    ����    IU    ����    ����    ����    �W    ����    ����    ����    �\    ����    ����    �����_�_    ����    ����    ����    ��    ����    ����    ����    |�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    q�    ����    ����    ����    ��    ����    ����    ����    F�    ����    ����    ����    U�    ����    ����    ����    ��    ����    ����    ����    >�    ����    ����    ����    ��    ����    ����    ����    {�    ����    ����    ����    ��    ����    ����    ����    <    ����    ����    ����    �	    ����    ����    ����    �        �        ����    ����    ����    <"    ����    ����    ����    B    ����    ����    ����    �I����    	J        ����    ����    ����    �L����    eM        ����    ����    ����    �S    ����    ����    ����tjzj    ����    ����    ����6k<k    ����    ����    ����    ��    ����    ����    ����    >�    ����P."�   ��                           ����    ����    ����    �    ����    ����    ����    %�    ����    ����    ����    Ƽ    ����    ����    ����    b�    ����    ����    ����    @�    ����    ����    ����    k�    ����    ����    ����    P�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    D�    ����    ����    ����    H�    ����    ����    ����    ��    ����    ����    ����    ��        e�        ����    |��    ����            z        ����    ����    ����    n    ����    ����    ����    	    ����    ����    ����    �    ����    ����    ����� �     ����    ����    ����    �&    ����    ����    ����    �:        �9        ����    ����    ����    CA    ����    ����    ����    �B    ����    ����    ����    �E    ����    ����    ����    oH    ����    ����    ����    �Y    ����    ����    ����    �o    ����    ����    ����    ;r    ����    ����    ����    �    ����    ����    ������    ����    ����    ����]c    �����."�   �                           ����    ����    ����     w    ����    ����    ����    ly    ����    ����    ����    T|    ����    ����    ����    ��    ����    ����    ����    b�����    ͊        ����    ����    ����    "�����    Y�        ����    ����    ����    �        �        ԑ            ����    ����    ����    �    ����    x���    ����    ��    ����    x���    ����    C�    �����."�   Ȫ                           ����    ����    ����    ��	    ����    ����    ����    ��	    ����    ����    ����    ��	    ����    ����    ����    
�	    �����."�   x�                               ��    ��       ̫�        p�    ����       y�        ��    ����       u�        ����    ����    ����    �N
    �N
�N
        ����    ����    ����    8R
    9Q
FQ
        ����    ����    ����fV
lV
    ����    ����    ����X
X
    ����    ����    ����Y
Y
    ����    ����    �����`
�`
    ����    ����    ����_a
la
    ����    ����    �����a
	b
    ����    ����    �����b
�b
    @           >d
����    ����                  P�"�   `�   p�                       ����P/"�   ��                           ����    ����    ����    ��
    ����    ����    ����G�
w�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���R    �          ذ ܰ � �� �   AnimaWrapper.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T            �     
  $  m  �  J    #   ̤    .?AVBaseData@@         N�@���D        u�  s�          ̤    .?AVtype_info@@          �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                             �   ����   ��������    �����
                                                                                  `�P�    ��������                       ��������������������                                                                                                                                                                                                                                                                                                                                            abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     `��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            ����C   ���� �������������������������������������������t�h�`�X���P�H�@�4�(�����������	         ��������������t�d�P�8� ������������������������t�h�T�<�,��������������������p�@�(�                                                                                                                                                                   ��            ��            ��            ��            ��                              8�         >�BD��                                            @�@�`�                �p     ����    PST                                                             PDT                                                             p���                                ����        ����                                                                                                                                                                                                                                                                                                                                                                     Q�����         ������������                    �                                                                                                                                                                                                                                                                     �                            .   .   0�������������������4���������������8�                     >@    ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                      @          ���5      @   �  �   ����                         ̤    .?AVbad_exception@std@@         ̤    .?AVexception@std@@                .          ����                   �D        � 0                          �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                            ̤    .?AVbad_cast@std@@      ̤    .?AVbad_typeid@std@@        ̤    .?AV__non_rtti_object@std@@                                                                                                                                                                                                                                                                                                                                         <         � L          � (                     \ n � � � � � � � 
  . @ Z r � � � � � �  " 2 B P b r � � � � � � �   $ < L d x � � � � � �   , B T ` p � � � � � � � �   2 J V d p � � � � � � � �   * < L \ n � � � � �                                                                                                                     � �                                             \ n � � � � � � � 
  . @ Z r � � � � � �  " 2 B P b r � � � � � � �   $ < L d x � � � � � �   , B T ` p � � � � � � � �   2 J V d p � � � � � � � �   * < L \ n � � � � �                                                                                                                     � �                                             =LoadLibraryExA  GetModuleFileNameA  EGetProcAddress   IsDebuggerPresent KERNEL32.dll  MessageBoxA  GetActiveWindow USER32.dll  �GetCurrentThreadId  � DecodePointer �GetCommandLineA �GetTimeFormatA  �GetDateFormatA  yGetSystemTimeAsFileTime � EnterCriticalSection  9LeaveCriticalSection  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter � EncodePointer GetModuleFileNameW  �HeapValidate  �IsBadReadPtr  GetLastError  R CloseHandle oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection RtlUnwind �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  �InterlockedIncrement  sSetLastError  �InterlockedDecrement  �GetCurrentThread  ExitProcess aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId gMultiByteToWideChar �RaiseException  MlstrlenA  ?LoadLibraryW  IsProcessorFeaturePresent hGetACP  7GetOEMCP  rGetCPInfo 
IsValidCodePage �GetTimeZoneInformation   FatalAppExitA %WriteFile �OutputDebugStringA  $WriteConsoleW �OutputDebugStringW  -SetConsoleCtrlHandler �HeapAlloc �HeapReAlloc �HeapSize  �HeapQueryInformation  �HeapFree  �SetStdHandle  WFlushFileBuffers  �GetConsoleCP  �GetConsoleMode  �ReadFile  � CreateFileA bFreeLibrary �InterlockedExchange GetLocaleInfoW  JGetProcessHeap  �VirtualQuery  -LCMapStringW  iGetStringTypeW  fSetFilePointer  SSetEndOfFile  GetLocaleInfoA  IsValidLocale EnumSystemLocalesA  �GetUserDefaultLCID  � CreateFileW d CompareStringW  VSetEnvironmentVariableA                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                 0  �              	  H   X  Z  �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel>
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPAD   p   P2V2z2�2�2�2�2�23%3:3?3E3L3Q3�3�3�3
444:4@4V4[4e4k4p4x4�495>5E5�56|6�6Z7�7p8�8�8�9l:�:;;�<$>H>T>�?  H   /1�12�2�2h3�3w45�5�5�67�78�89�9:�:�:k;�;K<�<+=�=>�>?�?     T   C0�0+1�122�2+3�344�4�5
6�6;7�7�7�=�=�=�=�=%>0>K>P>Y>^>c>�>�>x?}?�?�?�?�?�? 0     �34�4/5�5"6@;h;t;�;k<�< @ h   �1�1�1383D3�3�3�3�3�3�3�3/4�4�4�4�4�5�5�5�5�5�5�56�6�6�6�67�7o8�8o9�9?:�:�:�;_<�<b=�=e>�>?�? P ,   0�0�0o1�1n2�2�3K5r5�9::<,<8<L>�? ` T   10T0`0�0�0 1�1�1�1=2�2"3�3s4�4#5E5�5�5{6�6�7�7d8�8R9�9r:;+<�<=�=>�>?�?   p T   0�0�0�01o1�1o2�2o3�3F4�4/5�5.6�67�78�89�9�9d:�:K;�;+<�<={=�=[>�>;?�?   � D   �6�6*7P7\7h788!8&8W8b89�9::�:�:�:�;�;><d<p<�<b=l>�>L?�? � L   +0�01�12�2�2X3�3�4�4T5�5D6�6R7�7b8�8T9�94:�:;�;�;~<=}=�=Z>�>:?�? � L   0�0�0)2L2X2�2J3�3B4�4-5�5)6�6*7:7=8-9�9:}:�:F;�;D<�<+=�=>{>�>[?�? � P   ;0�01�1�1k2�2K3�3+4�45{5�5_6�6O7�7K8�8r9�9|:�:\;�;;<�<=�=>�>?�?�?   � P   k0�0K1�1+2�23{3�3k4�4[5�5W6�6D7�7+8�89�9�9t:�:T;�;;<�<2=�=J>�>�> ?�?   � P   ?0�01�12�2334�4"5�5'6�627�7/8�8*9�9
:v:�:n;�;!<D<P<�<
=o=�==>�>?�? � `   0�0�0k1�1V2�2�23<3H3�3�34�4G5�5&6�6�6f7�7/8�89o9�9J:�:-;�;<�<�<r=�=�=�=:>�>)?�?�?   � h   j0�0M1�12T2x2�2�2F3�3j4�4m5�5M6�6-7�7
8z8�8V9�9G:q:�:�:�:�:7;a;�;�;�;�;'<Q<t<�<�<�<=�=S>??�?     L   K0�0K1�1/2�23�3�3O4�4&5�56�667�7M8@9d9p9�9J:�:0;�;M<�<F=�=B>�>[?�?  d   �0�0$1*1P1�1�1.232<2A2F2w2�2)3�3�4�4�4O586\6h6�6�7�7�7�8�8�8�9�9�9O:�:J;�;<�<=�=�=m>�>M?�?   l   &0�0
1v1�1O2�2"3�3�3f4�4$505�56}6F7�7�78r8C9�9�9�9:D:P:\:h:�;�;�;�;�;<%<�<�<�<=q=�=�=>4>@>B?�? 0 H   h0�01$1�1�1n23z3�3O4�4*5�5�5j6�6a7�7�7�7]8�8�9�:�:;k<�<�=?�? @ t   0�0�14A4J4�4&535�5�5�5666�6�6f7�7�78.:4:::@:F:L:�:�:�:�:�:;;;<<5<:<?<�>�>?W?`?�?�?�?�?�?�?�?�?   P �   0&0P0U0Z0�0�01 1T1]1�1�1�1h3m33�3�3�3�3�344I4N4S4x4�4�4�4�45)656b6g6l6�6�6�6%7.7X7]7b7i9t9�9�9�9�9b;�;�;�;�;�;�;V<^<o<x<�<�<�<�<== =:=h>m>>�>�>�>Y?l?�?�?   ` �   �2�2 3�3444444%4)4/43494=4C4G4M4Q4W4[4a4e4�4�4�4�4z6�6�6�6�6�6�6�6	7/7M7T7X7\7`7d7h7l7p7�7�7�7�7�728=8X8_8d8h8l8�8�8�8�8�8�8�8 9999V9\9`9d9h9;e;j;o;�;�;�;9=J=b=s=�>Y?^?c?�?�?�?   p �   ,2�2�2�2333�3�3�3�3�3�3Z4_4d4�4�4�4 5%5*5�5�5�5�5�5�5t8�8�8�8�8�8�8&9+909l9x9�9�9�9::F:s:x:}:M;Y;$<0<]<b<g<�=�=&>2>_>d>i>�>�>???u?�?�?�?�? � �   0)0V0[0`0�1�122"2�2�2�2�2�2-393f3k3p3�3�3+40454�4�4�4�4�4F5R55�5�5�5�5&6+606�6�6�6�6 7l7x7�7�7�788F8K8P8�8�8�8�8 9l9x9�9�9�9�:�:�:;;�;�;�;�;�;{<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ===   � l   �344�5�5�5!6�67�7�7v8�8�9�9�:�:(;,;0;4;8;<;@;D;H;L;P;�;�;�;�;�;�;�;�;R>^>�>�>�>??B?K?u?z??�?   � �   00&0+000N0S0X0^5/686b6g6l6�6�6�6�6�6�8.:�;�;�;�;�;�;�;<<<(<2<@<F<v<<�<�<�<�<m=~=�=�=�=�=G>h>q>�>�>?)?G?T?�?�?�?   � �   �0�01�1�1�1�1�12�23�3�3�3�34�4�4�4�4�4E5u5�5�5�5�5�56#6(6O6X6�6�6�6�6A7Z7c7�7�7�788J8S8\8�8:P:`:e:j:o:�:�:�:�:[;g;�;�;�;�;�;�;�;<<.<:<f<�<�<�<�<==9=>=C=v={=�=�=�=�? � �   �0�0�0�01c2�3�3�334;4D4T4`4v4�4�4�4�4�4�4�4�45595T5�5�5�56_6j6s6{6�6�6�6�6�6�6�6�6�6�67727Q7F9X:]:o:o;x;�;�;�;�;�;�;�;�;�;�;<)<F<K<�<�<==$=E=e=�=�=�=>C>Q>�>�>�>�>�>????+?4?:?C?H?N?V?\?�?�?�?�?   � �   @0J0V0r0�0�0�0�0�0�0�0�0�0�3�3�3�3�34#4(455/5�5�5�5�5�5�566*6J6v6�6�6�6�6�607<7R7d7�7�7�7�78n8t8�8�8�8�89\9h9�9�9�9�9�9�9�9:::3:D:w:�;�;<5<A<n<s<x<�<�<�<�<�<�<�<�<==i=u=W>c>�>�>�>??�?�?�?   � �   80=0O0c0�0�0�0�0�0110151R1W1�1�1�1�1A2p2�2�23F3}3�3�3!4x4|4�4�4�5�5�5�566D6I6N6[6t6�6�6�6�6H7M7_7�7�7�7�7�7�7�79989=9O9):G;S;v;�;�;�;�;�;�;<<.<k<=7=[=f=C>O>|>�>�>�>�>�>�>�>?!?N?S?X?�?   � �   11/1[1`1�1�12*2U2w2�2�2�23A3�3�3�3�4�5666N6�67,717�7�7�7�7�7898]88^:j:�:�:�:�:�:;;";�;)=F=w=�=�=�=�=>>E>Q>~>�>�>\?   �   �1�1�12w2�2�2�2>3J3w3|3�3X4]4o4�4�4�4555B5Z5c5�5�5�5�5667'7]7p7�7	88<8A8F8�8�889=9O9x;};�;�;�;�;<3<O<y<�<�<�=�=�=�=�=2?>?    �   n0x0�0�0�0�1�1�1�1�1�1�1�2�2�2C3�3�34^4e4�5�5�5�5�56Y6|6�6�6�6�6�6p7y7�7�7�7
88�9�9�9�9�9<:m:y:�:�:�:;;G;L;Q;�;�;�;1<=<j<o<t<�<�<�<�<�<*=3=�=�=�=�=�=�=�=�=�=�=�=�=�=     �   000a0o0�0�0�0�0
1(1?1W1q1~1�1�1�1�1�13!3,4�4�465>5]5g5�5�5s667�7�7�7�7�7V8h8�8�899>9C9H9�9�9�9�9�9t:�:�:I;U;�;�;�;9<@<N=U=�>�>g? 0 h   20�0?1K1{1�1�1`2�2�233H3O3�8�8�8�8�8�8�8�8�8�8�8 999 9$9(9,909d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9 @ `  (1-1?1p1y1�1�1�1�2�2�2 3P3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444(4-434=4G4S4_4d4v4{4�4�4�4�4	5'5K5R5v5�5�5�5�5�5�5�5�56696C6H6M6W6\6a6k6p6u66�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6777#7*7/757<7A7F7M7R7l7r7y7�7�7�7�7�7�7�7�8�8�8�8�8�8�8�8�89993999F9�9�9�9z:�:�:�:�:�:�:;�;�;�;�<�<�<4==='>5><>F>M>T>`>g>n>>�>�>�>�>�>�>???3?@?E?S?[?s?   P �   g0�0�0�0�0�011'1.1=1G1U1Z1a1k1o1y1�1�1�1�1222@2M2Y2i2p2�2�2�23333Q3V3c3h3v3�3�3y44�4�4�4K6W6�6�6�6�6�6�6�6�6�67{7�7�7�7�7�7�7�7 8%8*8B8�8�8�89!929v9�9�9�9�9�9�9::�:�:�:�:�:�:�:�:;U;�;�;	<   ` �   q0�0�01*1M1�1�1�1�1�1�122#2V2]2c2�2�2�2�2�2�2�2�233(343D3�3�3�4�4�4�6�67727|7�7868q8�8�8 919Y9::/:n:�:�:�:0;�;�;�;,<`<e<�<�<=
===#=>=D=M=V=[=f=�=�=�=�=�=�=�>�>�>�>2?l?�?�? p �   00S0Z0y00�0�0�0�0�0�0�011F1V1Y2^2z22�2)6t6�6�6�6�6�6�6777~8�8�8�8�8�8�8,91969x9�9�9�9�9�:�:�:�:�;�=�=�=�=�=�=>0>5>:>v>�>�>�>�>   � H   �6D7P7}7�7�7�7�7�7�7�739?9l9q9v9�9�9�9�9�9)<x<�<�<�<�<�<�<==#= � �   �0�0�0Q2Z2�2�2�2�2�233I3N3S3�3�3414:4d4i4n4�4�4�5�5�5�5$666A6Y6b6o6777s7�7�7	88D8O8[8�8�8�8�8�8999"9,9T9H:W:�:�:�:�:�:�:�;�;G<�<	=K=e=�>�?�?   � �   00000�01l1�166<6X6t6�6�6�6�6/7G7�7�7�7
8&8O8u8�8�8?9�:�:;�;=h=m==�=�=�>�>�>�>�>�>�>�>???]?d?h?l?p?t?x?|?�?�?�?�?�?�? � �   B0M0h0o0t0x0|0�0�0�0 11111111f1l1p1t1x1Y7b7�7�7�7�7�78,81868M8�8�8�8�8�8�8]9f9�9�9�9�9�9:::K:T:~:�:�:�:�:v;�;�;�;�;�;�;�;�;<<x<}<�<===}=�=�=�=�=�=�=�=�= >
>>>>B>L>[>d>j>y>�>�>�>�>�>�>�>�> ?3???p?y?�?�?�?�?�?�?�?   � �    000�0�0�1�1�1�3�3�3�4�4�4�4�4�4�45
555$5,545Q5Y5a5i5q5}5�5�5�5�5�5�5�5�5�5�56
666�6�6�6�677+797Q7_7�7�7�799�9�9U:d:�:�:�:�:�:�:�:�:;;;';-;6;>;J;V;[;c;l;W<`<�<�<�<�<�<�<==�>�>?+?0?5?^?g?�?�?�?   � P   I0R0|0�0�0�0�0�0�0�033X7a7�7�7�7�7�78	8899�:<(<�=�=&>2>�?�?�?�?�? � �   %0.0�0�0�011�1�1�1�2�2�223<3�3�3L4Q4�4�4�45�5�5�5�6�6�6H8M8_8�8�8�8�8�8
99*9�9�9::%:3:�:�:�:�:�:�:
;;$;h;m;;�;�;�;</<b<=2=9=[=b=}=�=>>H>M>R>�>�>�>�>�>�>�>?�?�?�?�?�?   � $  00$0.0>0H0W0�0�0�0�0�01�1�1�1�1�12!2<2I2N2T2a2f2l2�2�2�2(3-32373j3v3�3�3�3�3�3�3�34444C4H4M4R4�4�4�4�4#5(5-525]5b5g5�5�5�5666696B6t6�67�7�7�788%878A8_8d8i8�8�8;;6;<	<<"<'<O<U<p<}<�<�<�<�<�<===R=W=\=a=�=�=�=�=�=�=�=�=$>5>:>?>D>m>r>w>|>�>???M?R?W?\?�?�?�?�?�?�?   �   0!0&0+0N0W0�0 1�1�1�1 222S2Z2i2�2�2�233J3Q3[3m3w3�3�3�344�6�6�6�6�6�6�6b7l7r7}7�7�7�7�7�7�7�7�7�7	88880858=8D8W8\8�8�8�8�8�8W9�9�9�9�9�9�9:,:0:4:8:<:X:\:h;m;;�;�;�;�;�<�<�<�<�<�<
='=D=�=�=�=�= >>�>�>�>\?`?d?h?l?p?    �   r0�0�0�091h1t1z1�1�1�1�1�1�1�1�1�1�1�1�1�1�1
2222'2.23292D2N2U2^2e2�2�2�2�2�2�2334+4X4]4b4�4�4�4�4�499;9@9E9�9�9�9�9�9�9�9&:+:0:A;J;t;y;~;�;�;
<<=<B<G<�<�<=*=3=]=b=g=�=�=   �   00/0H0y1�1�1�1�1�1�162=2W2^2�2X3�3�3�3�3�34$4N4S4X44�4�4�4�4�4q5�5�5�56%636?6z6�6�6�6@8~8�8�8�8�8�8�8 99�9�9�9�9�9�9�9:":.:I:Y:e:�:�:�:�:�:0;6;d;i;n;�;�;�;�;�;L=U==�=�=�=�=�=�=>�>�>E?L?x?�?�? 0 �   >0E0T0�0�01(1R1W1\1�1�1�1�1�1s5|5�5�588X8]8o8�8�89U9�9�9�9:5:;:D:Y:�:�;�;�;<$<2<H<�<�<==8=D=P=f=>*>6>n>s>x>�>�>�>�>�>?'?�?�?�? @ �   0 0�0�0�0
1&1[1y1X2]2o2�2�2"3-3�3�3�3�3�3&4I4R4|4�4�4�4�4�4�4�45:5W5a5�5�5x6}6�6�6�6�62777<7b7z7�7�7�7�7�7D8M809t9}9�9�9�9�9::T:Y:^:�:�:;;6;�;�;�;�;�;<�<�<e=�=�=�=>>:>�>�>�>   P �   00H0d1n1�1�2�233:3�3�3�3487=7O7�7�7�7�7�7�7"8:8C8x8}8�8�8�8�8�8�8*9s9|9�:�:�:;!;&;L;d;p;�;�;�;�;�;<"<'<Z<�<�<�<�<�<�<3=?=w=|=�=�=>=>I>�>�>�>�>�>?R?y?�?�?   ` |   0+0e0�0�0�0'1l1�1�1�12(2F2&303:3s3�3u4�4�45I5w5�5�5 6X6v6�6�6�67278'818o8�8�89�=�=�=�=�=�>�>�>�>�>?"?'?�?�?   p �   x0}0�0�0�0�0�0�011=1j1o1t1�1�1�1�1�1]22�3�3�3�4�4�4�4�455�5�5�5�5�5�6�6�677078i8�8�8�8�899:9h9�9�9�9%:F:g:�;�;!=�=�>�>I?U?   � h   �0�0(1P11�1�12252W2�2�2�2�2�2�2�2034383<3@3D3H3L3P3T3�8�8�8�8�899C9H9M9�>�>�>�>�>�>?2?7?<? � �   �1a2m2�2�23�3�3�3444-4�4�4�4�4�4�5�5�5�5�5S6v6�6�6�6�6�6:}:�:�:�:�:F;X;�;�;�;�;.<3<8<z<�<�<�<�<d=�=�=�=">'>,>w>�>�>$?)?.?�?�?   � |   �0�0(2/23�374�4�455$5�5�6�6�6�6�6�6�<�<�<�<�< =$=(=,=0=4=8=<=@=D=H=L=P=T=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= � L   L829>9n9s9x9�9:R:d:�:�:�:�:�:5;A;q;v;{;�<�<>$>T>Y>^> ??<?A?F?�?   � �   40@0p0u0z0E1L1]2i2�2�2�2�3�3�3�3�3A5M5}5�5�5x6�6�6�6�6�7�7�8�8�9�9�9�9�9�:�:�:�:�:�;�;(<-<2<�<=8===B=&>2>b>g>l>6?B?r?w?|?�? � �   &121b1g1l162B2r2w2|2�2i3+474g4l4q4;5G5w5|5�56(6X6]6b6N7Z7�7�7�7Q8]8�8�8�8<9�9:6:;:@:v:�:;;F;M;�;�;==@=E=J=> >P>U>Z>8?D?t?y?~? � p   H0T0�0�0�0{1�1�1�1�1�2�2�2�2�2�3�3�3�3�3�4�4�4�4�4�5�566!6�6�6'7,71788=8B8G899M9R9W9�>�>�>�>�>�?   � h   �0�011 1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222 2$2(2,2024282<2@2D2H2�2�2�2�2�2�2�2�2     �   x3}3�34 4)404�4�455)5A5F5�56666t6�6�67�7�7R8n8y8�8�8�8�8�8�8�8999m9r9w9~9�9�9�9�9�9�9�9�9:":':;;!;8;=;O;<<<6<=<�<�<�<�<=.=3=8=b=h=�=�=�=�=�=�=�=&>/>K>f>k>p>~>�>�>�>�>|?�?  x   #0�0�0�0�0\1w1�12	387G7W8t8�8�8�8�8�8�89U9#:*:�:�:�;�;�;�;�;�;�;�<�<�<	==1=?=X=n=�=�='>-><>E>N>W>a>u>?e??     ,   m0v0�0�0�0�1�2�3�4w5W677'89:�:�>I? 0 X   �0)2�3�3�3�3�34%4O4T4Y4�4�4�4�4�4�45-52575�6H7M7R7y9�9�9�9�9�9�9:8;�<�<�=�=�= @ (   C2�2�2A3�3�3$46�6�627�7�7�7�7�7 P    �?   ` h   0c0�1�1�1�1�12!262B2n2W4u4�4�4�4W55�509�9�9�9�9%:�<�<�<�<=3=R=q=�=�=�=�=>�>�>�>�>?,?�?�?   p �   J1S1}1�1�1�1�1,242q2z2�2�2�23&3�3�3�3'404Z4_4d4�4�4�5�5656>6h6m6r6�6�6�6�6�6�7�7�7�7w8�8999�9�9:	::b:n:�:�:�:;;!;�;�;�;�<�<�<�<�<?=K=x=}=�=	>>>�>F?\?w?�?�?   � x   20Z2t2�3�3�3"404>4�56�6�6�67^7l7�7�7�718\8h8�8�8�8�8�8�8�899/9D9H9`9e9r9�9�9�9/:=:�:�;�;)<�<h>m>>�>G?�?�?�? � `   90E0r0w0|0�0I1_1�1�1�2�2�2�2�23,3�3]4y4�4�4�4�48�8f9k9p91;�;<r<�<�<�>?(?M?R?W?\?�?�? � �   0/0�0�0�0
1<2�2�2�2�24)4.434�4�4�4�5�5�5z66�6�67 7%7j7o7t7�7�7�7�8�8�8�8*9�9�9�92:U:^:�:�:�:�:�:�:;!;&;b;�;�;�<�<=%=X=v=�=�=�=;>k>�?�?�?�? �   ,0�0�0�0�0�0�0�01111%1}1�1�1�1�1�1�1�12"22�2�2�2�2�2�2�2�2�23�3,494b4l4�4�4�4�4�4�4�4�4�45d5u5�5�5�5�5#6�6�6�6�6�61768D8h8q8�8�8�8�89!9F9O9X9c9l9q9�9�9�9�9�9�9�9�9�9�94:S:`:�:�:�:�:�:;";5;:<I<R<x<<�<�<=+=3=9=]=o=�=�=�=�=>>%>K>R>X>a>y>�>�>�>�>�>�>)?4?K?V?�?�?�?   �   040B0Q0Z0�0�1�1�1�122#2H2P2i2�2�2�2�2333)343C3i3v3~3�34@4D4H4L4P4T4X4�4�4�4�4�4�4�4�4�4�4�4�4�4P5T5X5\5`5d5h5�7�7�78	88.878Y8e8s8|8�8�8�8�8�889I9\9g9�9�9�9�9�9':.:4:C:Q:Y:�:�:�:�:�:$;5;P;c;p;y;<_<�<�<�<�<�<�=>>>�>�>�>�>�>�>�>?? ?K?^?g?�?�?�?�?   � �   050=0H0P0X0�1222,252N2\2o2|2�2�2�2�2�2�2,3:3[3d3j3r3{3�3�3�3�3�3�354�4�4�4�4�4�4Y5s5�5�5�5�5�5�5	66'6/646G6T6c6l6�6�6�6�67*7l7z7�7�7|8�8�8�8�8�8�8�8�8�8$9U:�:�:�:�:�;7<@<p<t<x<|<�<�<�<�<�<�<�<�<�<�< � $   �1�1�56|7!8G8T8{:�;a<=D>V? � x   	1�1w2"3�3�3�9�9�9�9�9�9�9:O;�;<<<3<:<�<�<�<�<�<�<�<�< ===!='=5=B=K=T=�=�=�=�=�=�=�=�=>)>�?�?�?�?�?�?�?    	 �   0]2k2t2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2@3D3H3L3P3�3�3�3�3�3�3�3�3�3|6�6�6�6�6�6�7�7�7�7�7�7�7*8�8�8�8�8 9'9�9�9�9 :::::�:�:�:�:2;;;L;g;~;�;�;Q<k<r<�<�<�<�<�<=G=P=U=o=v=|=�=�=�=�=�=�=>J>S>Z>�>�>�>�>�> ?????X?\?`?d?h?l?p?t?x?   	 <  �0�0�0�011'1,1]1�1�1�1�1�1�1�2�2�2�2�233)3G3U3h334&444=4m4�4�4
555U5\5a5s5�5�5�5�5�5�5�566&676I6[6m66�6�6�6�6�6787A7R7a7p7x7�7�7�78B8I8R8�8 959L9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::h:l:p:t:�:�:Z<e<m<�<�<�<�<�<�<�<�<�<�<=t=x=|=�=�=�=�=�=�>�>�>�>�>�>?#?/?8?W?^?g?�?�?�?�?�?�?�?�?�?�?  	 �   <0c0p0~0�0�0�0�0�0�0�0i1�1�1�1�12M3�5�5�5�5Q7Y7_7�7�7�7�7�7�78888'8_8n88�8�8�8�899#9::^:g:�;�;�;B<K<s<�<�<\=z=�=�=>>!>�>�>   0	 �   �2�2�2�2�23-3:3B33�3L4�4�4�5[7�7�7�8�8�8�8v9�9�9�9:F:S:[:m:z:�:�:�:�:�;<2<@<I<�<F=f=�=�=�=�=>&>F>f>�>�>�>�>?"?F?n?�?   @	    �3:):�; P	    �2D56�6+8�<?r? `	 X   �0�1�1�2�2h4�576e6�6�6�6�6�6�6�6�67.757�7Y:b:�:�:�:Z;�;r<=w>>? ?M?R?W?�?�?   p	 �   0"0O0T0Y0�0�0h1p1�1�1�1�1�1�3�3�3�3�344V4_4�4�4�45585a5j5�5�5�566F6o6x6�6�6�6�6�6o8x8�8�8�8�8�89!9&9�:;r;~;�;�;�;�;�;+<0<5<^<�<�<�<�<(=-=2=p=w=�>�>�>�>�>B?N?{?�?�?�?   �	 �   00{0�0�0B1N1{1�1�1�1�1K3�3{4�4�4�4�4�4�4555S5[5�5�5�5�5�56#6M6R6W6!7-7Z7_7d7�9�9�9�9�9	::B:G:L:�:�:�:�:	;;;R;^;�;�;�;�<�<�<�<�<Y>�>�>�>�>�>�?   �	 �   �0�0'1�2�5�5�5�5�566�6�6�6�6�6)717�7�7�7 8-82878�9�9�9�9�9#:+:j:s:�:�:�:;$;Q;z;�;�;�;�;1<8<e<�<�<�<�<�<==�>�>�>�>�>??H?M?R?   �	 �   [1�1"2.2[2`2e2�2�2�2�2�23H3O3�3�3�3�3�3#4+4Y5e5�5�5�5�5�5+60656w6�6�617�7�7�7
878<8A8�8�8:}:K;T;~;�;�;�;�;�;�;�;%<-<r<{<�<�<�<�<�<!=&=+=�=
>7><>A> �	 �   �0�0�0�0�0�012171<1w11�1�1�122F2R22�2�2�3�3�3�3�3l5�5�566#6e6q6�6�6�6Q7�7�7A8H8W9^9�:�:v;?<�<r=~=�=�=�=�>??F?M?{?�? �	 l   5555555 5$5(5,5054585P5T5X5\5`5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5/<;<h<m<r<�<�<�<�<�<�>?8?=?B?�? �	 �   0@0r0�0�0�0�0�0�0111'1.13181B1I1N1S1]1j1o1u1}1�1�1�1�1�1�1�1�1�12*212K2V2]2u2|23�3�3�3�3�3�344 4�5�5�5�5�5�6�6�6"7H7M7_7�78"8)8�8�8�93:8;=;O;�;�;�;�;�;�;<3<<<q<v<{<�<�<�<�<=?=k=t=??   �	 �   +0200�0�1�1�1A2d2m2�2�2�2�2�2�2(3-323k3�3�3�4�4�45:5X5�5�5�56%6O6T6Y6�6�6�6�6�6�67/787b7g7l7�7�7�7�89�9�9�9�9�9:9:Z:t:�:�:�:�:	;<<I<N<S<k<q<�<�<===#=�=�=�=�=�=�=�='>,>1>g>p>�>�>�>   �	 �   *0H0T0�0�0�0�0�0�0�0�0 1,1Y1^1c12-2x2�2�2�2�233a3j3�3�3�3�8�8{9�9�9�9�9�9�9�9I:�:�:�:�:�:(;0;�;�;�;�;<<<�<�<==E=r=�=�=�=�=�=> >~?�?�?  
 h   0�011Y1|122D2I2N2v4~4�4�4575@5j5o5t5�7�7�8�8�9�9E:M:�:�:;;s;{;�;�;�;�;�;:<F<s<x<}<�>�>�?   
    �0�0�0M1w1|1�1v;�;    
 T   �3�3�4q5}5�5�5�5F6q7x7�8�8�9�9�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>???X?\?`?   0
 4   Y2c2�2i3i9�91;6;;;@;�;�;�;�;�;�;�;�;,<1<6<;< @
    05=5j9�9
:�=�=�= P
     h0m00(4-4?487=7O7�8�8�8 `
 h   x0}0�011/1�1�1�1X2]2o2�34]4�4�6�6�6	7M7V7�7�7�7�7�7 8%8*8�=�=�>�>�>�>�>'?0?Z?_?d?�?�?�?�?�?   p
 `   �1�1�1�1�355555�7�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==   �
 D   �0R1 2:2�2�2�2�2�2�2�4�4|5�546�7;;l;�;�=�=�=>?g?�?�?�?�? �
 l   c0�0W2^2�2�2�2�2�2�23}3�3�3�3�344A4F4K4�4)5s55�5�5�56�6�6�7�7�8�8�9�:;�;�;�;<<�<f=m=�=�=�=�= �
 l   h3t3�3�3�3�3 44444444 4$4(4,404H4L4P4T4X4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4L>2?>?n?s?x?�?�?�?�?   �
 p   0L1�1�2�2�2�2�2�3�3�3�3�34�4�466I6N6S6F7R7�7�7�7�8�8/94999,:8:h:m:r:6;=;�<�<9=E=u=z==K>W>�>�>�>�?�? �
 �   0"0'0�0�0/14191�1�2�23!3&3�3�3.43484�4J56$6T6Y6^6*767f7k7p788G8L8Q8>9J9z99�9C:O::�:�:.;�;�;'<,<1<g<s<�<=9=@=w=~=�>?7?<?A?   �
 x   00I0N0S021>1n1s1x1D2P2�2�2�2w3�3�3�3�3�4�4�4�4�4�5�5�5�5�5�6�6�6�6�6�7�788!8�8�8)9.939::?:D:I:;!;Q;V;[;   �
 p   �0�0�0�0�0�1�2�2�2�2�2X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4\4`4d4h4l4p4t4 �
 X   �3�3�34484=4B4	5j5v5�5�5�6�6�8�8�89999B:W:l:�:�:�:�:;,;|;�;(<h<�<i=�?�?     �   0�0�0.1�1"2*3�3�3�3j4�4�4:5^5�5�6�6�6�7z8�8"9D9;;7;<;A;w;�;�;�;�;�;�;<"<'<�=>#>M>R>W>�>�>�>�>!?'?/?=?C?V?�?�?�?�?�?�?�?�?�?  `   00%010�0�0�0M1]1�1�1222q24a4q4�4A5j5o5t5i6r6�6�6�6�6�67 7%7o;x;�<�<|=�=? ?J?O?T?   �   �5�5 666666$6*60666<6B6H6N6T6Z6`6f6l6r6x6~6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677777 7&7,72787>7D7J7P7V7\7b7h7n7t7z7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7j>�>�>�>�>
?2?j? 0    �?�?�?�? @ �   0060p0v0�0�0�0�00161p1v1�1�1�1�10262p2v2�2�2�2�20363p3v3�3�3�3�30464p4v4�4�4�4�40565p5v5�5�5�5�50666p6v6�6�6�6�60767p7v7�7�7�7�70868p8v8�8�8�8�80969p9v9�9�9�9�90:6:p:v:�:�:�:�:0;6;p;v;�;�;�;�;0<6<p<v<�<�<�<�<0=6=p=v=�=4>�>�>�>�> ??@?F?�?�?�?�? P �    00@0F0�0�0�0�0 11@1F1�1�1�1�1 22@2F2�2�2�2�2 33@3F3�3�3�3�3 44@4F4�4�4�4�4 55@5F5�5�5�5�5 66@6F6�6�6�6�6 77@7F7�7�7�7�7 88@8F8 p �   1111111 1,1014181<1@1D1H1T1X1\1`1d1h1l1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222222$2(2,2024282<2@2L2P2T2X2\2`2d2h2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�5 66699$:   �    L:P: �    �2   �    �4�4<6@6D6`>d>h>l>p> �    �<�< �     �4�4�4�4�4�499999        �7�7�7     4   L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< @ ,   H<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<   ` �   000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6   p    �>�>�>�> � �   �5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 9999P<T<X<x<|<�<�<�<�<�<�<�< � h   T9X9l9t9|9�9�9�9�9�9�9�9:::$:(:0:H:T:l:�:�:�:�:�:�:�:�:�:�:�:;;,;4;8;@;X;p;t;�;�;�;�;�;�;   �    1 1@1`1�1�1�1�1�1 2 2@2`2�2�2�2�2 3 3@3`3�3�3�3�3�344@4L4p4�4�4�4�4�4�4�45@5`5�5�5�5�5 6 6@6`6�6�6�6�6�6�6 7@7`7|7�7�7�7�7�7808P8p8�8�8�8�8�8999(9`9�9�9�9�9�9::@:L:X:�:�:�:�:�:;0;P;p;|;�;�;�;�;�;�;�;�;<(<0<4<X<`<d<�<�<�<�<�<�<�<�<==$=(=D=H=\=�=�=�=�=�=�=>> � �   p0�0�0�0�5 66064686<6@6D6H6L6P6T6�:�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�>�>�>�>�>�>????D?H?L?�?�?   � D   �1�183<3@3D3H3L3P3T3X3\3h3l3p3t3x3|3�3�3�3�3�3(4p4�4P8p8�8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              